// Library - XB16TSMC65, Cell - ZFBAR4, View - schematic
// LAST TIME SAVED: May  8 15:13:02 2023
// NETLIST TIME: May 12 11:49:58 2023
`timescale 1ns / 1ns

module ZFBAR4 ( NR00, NR01, NR02, NR03, NR10, NR11, NR12, NR13, NR20,
     NR21, NR22, NR23, NR30, NR31, NR32, NR33, NR40, NR41, NR42, NR43,
     NR50, NR51, NR52, NR53, NR60, NR61, NR62, NR63, NR70, NR71, NR72,
     NR73, NR80, NR81, NR82, NR83, NR90, NR91, NR92, NR93, NR100,
     NR101, NR102, NR103, NR110, NR111, NR112, NR113, NR120, NR121,
     NR122, NR123, NR130, NR131, NR132, NR133, NR140, NR141, NR142,
     NR143, NR150, NR151, NR152, NR153, R00, R01, R02, R03, R10, R11,
     R12, R13, R20, R21, R22, R23, R30, R31, R32, R33, R40, R41, R42,
     R43, R50, R51, R52, R53, R60, R61, R62, R63, R70, R71, R72, R73,
     R80, R81, R82, R83, R90, R91, R92, R93, R100, R101, R102, R103,
     R110, R111, R112, R113, R120, R121, R122, R123, R130, R131, R132,
     R133, R140, R141, R142, R143, R150, R151, R152, R153, VDD, VSS,
     L00, L01, L02, L03, L10, L11, L12, L13, L20, L21, L22, L23, L30,
     L31, L32, L33, L40, L41, L42, L43, L50, L51, L52, L53, L60, L61,
     L62, L63, L70, L71, L72, L73, L80, L81, L82, L83, L90, L91, L92,
     L93, L100, L101, L102, L103, L110, L111, L112, L113, L120, L121,
     L122, L123, L130, L131, L132, L133, L140, L141, L142, L143, L150,
     L151, L152, L153, NL00, NL01, NL02, NL03, NL10, NL11, NL12, NL13,
     NL20, NL21, NL22, NL23, NL30, NL31, NL32, NL33, NL40, NL41, NL42,
     NL43, NL50, NL51, NL52, NL53, NL60, NL61, NL62, NL63, NL70, NL71,
     NL72, NL73, NL80, NL81, NL82, NL83, NL90, NL91, NL92, NL93, NL100,
     NL101, NL102, NL103, NL110, NL111, NL112, NL113, NL120, NL121,
     NL122, NL123, NL130, NL131, NL132, NL133, NL140, NL141, NL142,
     NL143, NL150, NL151, NL152, NL153, NRACK0, NRACK1, NRACK2, NRACK3,
     NRACK4, NRACK5, NRACK6, NRACK7, NRACK8, NRACK9, NRACK10, NRACK11,
     NRACK12, NRACK13, NRACK14, NRACK15, NVAL0, NVAL1, NVAL2, NVAL3,
     NX0, NX1, NX2, NX3, NX4, NX5, NX6, NX7, NX8, NX9, NX10, NX11,
     NX12, NX13, NX14, NX15, NX16, NX17, NX18, NX19, NX20, NX21, NX22,
     NX23, NX24, NX25, NX26, NX27, NX28, NX29, NX30, NX31, NX32, NX33,
     NX34, NX35, NX36, NX37, NX38, NX39, NX40, NX41, NX42, NX43, NX44,
     NX45, NX46, NX47, NX48, NX49, NX50, NX51, NX52, NX53, NX54, NX55,
     NX56, NX57, NX58, NX59, NX60, NX61, NX62, NX63, NX64, NX65, NX66,
     NX67, NX68, NX69, NX70, NX71, NX72, NX73, NX74, NX75, NX76, NX77,
     NX78, NX79, NX80, NX81, NX82, NX83, NX84, NX85, NX86, NX87, NX88,
     NX89, NX90, NX91, NX92, NX93, NX94, NX95, NX96, NX97, NX98, NX99,
     NX100, NX101, NX102, NX103, NX104, NX105, NX106, NX107, NX108,
     NX109, NX110, NX111, NX112, NX113, NX114, NX115, NX116, NX117,
     NX118, NX119, NX120, NX121, NX122, NX123, NX124, NX125, NX126,
     NX127, NX128, NX129, NX130, NX131, NX132, NX133, NX134, NX135,
     NX136, NX137, NX138, NX139, NX140, NX141, NX142, NX143, NX144,
     NX145, NX146, NX147, NX148, NX149, NX150, NX151, NX152, NX153,
     NX154, NX155, NX156, NX157, NX158, NX159, NX160, NX161, NX162,
     NX163, NX164, NX165, NX166, NX167, NX168, NX169, NX170, NX171,
     NX172, NX173, NX174, NX175, NX176, NX177, NX178, NX179, NX180,
     NX181, NX182, NX183, NX184, NX185, NX186, NX187, NX188, NX189,
     NX190, NX191, NX192, NX193, NX194, NX195, NX196, NX197, NX198,
     NX199, NX200, NX201, NX202, NX203, NX204, NX205, NX206, NX207,
     NX208, NX209, NX210, NX211, NX212, NX213, NX214, NX215, NX216,
     NX217, NX218, NX219, NX220, NX221, NX222, NX223, NX224, NX225,
     NX226, NX227, NX228, NX229, NX230, NX231, NX232, NX233, NX234,
     NX235, NX236, NX237, NX238, NX239, NX240, NX241, NX242, NX243,
     NX244, NX245, NX246, NX247, NX248, NX249, NX250, NX251, NX252,
     NX253, NX254, NX255, RACK0, RACK1, RACK2, RACK3, RACK4, RACK5,
     RACK6, RACK7, RACK8, RACK9, RACK10, RACK11, RACK12, RACK13,
     RACK14, RACK15, X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, X11,
     X12, X13, X14, X15, X16, X17, X18, X19, X20, X21, X22, X23, X24,
     X25, X26, X27, X28, X29, X30, X31, X32, X33, X34, X35, X36, X37,
     X38, X39, X40, X41, X42, X43, X44, X45, X46, X47, X48, X49, X50,
     X51, X52, X53, X54, X55, X56, X57, X58, X59, X60, X61, X62, X63,
     X64, X65, X66, X67, X68, X69, X70, X71, X72, X73, X74, X75, X76,
     X77, X78, X79, X80, X81, X82, X83, X84, X85, X86, X87, X88, X89,
     X90, X91, X92, X93, X94, X95, X96, X97, X98, X99, X100, X101,
     X102, X103, X104, X105, X106, X107, X108, X109, X110, X111, X112,
     X113, X114, X115, X116, X117, X118, X119, X120, X121, X122, X123,
     X124, X125, X126, X127, X128, X129, X130, X131, X132, X133, X134,
     X135, X136, X137, X138, X139, X140, X141, X142, X143, X144, X145,
     X146, X147, X148, X149, X150, X151, X152, X153, X154, X155, X156,
     X157, X158, X159, X160, X161, X162, X163, X164, X165, X166, X167,
     X168, X169, X170, X171, X172, X173, X174, X175, X176, X177, X178,
     X179, X180, X181, X182, X183, X184, X185, X186, X187, X188, X189,
     X190, X191, X192, X193, X194, X195, X196, X197, X198, X199, X200,
     X201, X202, X203, X204, X205, X206, X207, X208, X209, X210, X211,
     X212, X213, X214, X215, X216, X217, X218, X219, X220, X221, X222,
     X223, X224, X225, X226, X227, X228, X229, X230, X231, X232, X233,
     X234, X235, X236, X237, X238, X239, X240, X241, X242, X243, X244,
     X245, X246, X247, X248, X249, X250, X251, X252, X253, X254, X255
     );

inout  NR00, NR01, NR02, NR03, NR10, NR11, NR12, NR13, NR20, NR21,
     NR22, NR23, NR30, NR31, NR32, NR33, NR40, NR41, NR42, NR43, NR50,
     NR51, NR52, NR53, NR60, NR61, NR62, NR63, NR70, NR71, NR72, NR73,
     NR80, NR81, NR82, NR83, NR90, NR91, NR92, NR93, NR100, NR101,
     NR102, NR103, NR110, NR111, NR112, NR113, NR120, NR121, NR122,
     NR123, NR130, NR131, NR132, NR133, NR140, NR141, NR142, NR143,
     NR150, NR151, NR152, NR153, R00, R01, R02, R03, R10, R11, R12,
     R13, R20, R21, R22, R23, R30, R31, R32, R33, R40, R41, R42, R43,
     R50, R51, R52, R53, R60, R61, R62, R63, R70, R71, R72, R73, R80,
     R81, R82, R83, R90, R91, R92, R93, R100, R101, R102, R103, R110,
     R111, R112, R113, R120, R121, R122, R123, R130, R131, R132, R133,
     R140, R141, R142, R143, R150, R151, R152, R153, VDD, VSS;

input  L00, L01, L02, L03, L10, L11, L12, L13, L20, L21, L22, L23, L30,
     L31, L32, L33, L40, L41, L42, L43, L50, L51, L52, L53, L60, L61,
     L62, L63, L70, L71, L72, L73, L80, L81, L82, L83, L90, L91, L92,
     L93, L100, L101, L102, L103, L110, L111, L112, L113, L120, L121,
     L122, L123, L130, L131, L132, L133, L140, L141, L142, L143, L150,
     L151, L152, L153, NL00, NL01, NL02, NL03, NL10, NL11, NL12, NL13,
     NL20, NL21, NL22, NL23, NL30, NL31, NL32, NL33, NL40, NL41, NL42,
     NL43, NL50, NL51, NL52, NL53, NL60, NL61, NL62, NL63, NL70, NL71,
     NL72, NL73, NL80, NL81, NL82, NL83, NL90, NL91, NL92, NL93, NL100,
     NL101, NL102, NL103, NL110, NL111, NL112, NL113, NL120, NL121,
     NL122, NL123, NL130, NL131, NL132, NL133, NL140, NL141, NL142,
     NL143, NL150, NL151, NL152, NL153, NRACK0, NRACK1, NRACK2, NRACK3,
     NRACK4, NRACK5, NRACK6, NRACK7, NRACK8, NRACK9, NRACK10, NRACK11,
     NRACK12, NRACK13, NRACK14, NRACK15, NVAL0, NVAL1, NVAL2, NVAL3,
     NX0, NX1, NX2, NX3, NX4, NX5, NX6, NX7, NX8, NX9, NX10, NX11,
     NX12, NX13, NX14, NX15, NX16, NX17, NX18, NX19, NX20, NX21, NX22,
     NX23, NX24, NX25, NX26, NX27, NX28, NX29, NX30, NX31, NX32, NX33,
     NX34, NX35, NX36, NX37, NX38, NX39, NX40, NX41, NX42, NX43, NX44,
     NX45, NX46, NX47, NX48, NX49, NX50, NX51, NX52, NX53, NX54, NX55,
     NX56, NX57, NX58, NX59, NX60, NX61, NX62, NX63, NX64, NX65, NX66,
     NX67, NX68, NX69, NX70, NX71, NX72, NX73, NX74, NX75, NX76, NX77,
     NX78, NX79, NX80, NX81, NX82, NX83, NX84, NX85, NX86, NX87, NX88,
     NX89, NX90, NX91, NX92, NX93, NX94, NX95, NX96, NX97, NX98, NX99,
     NX100, NX101, NX102, NX103, NX104, NX105, NX106, NX107, NX108,
     NX109, NX110, NX111, NX112, NX113, NX114, NX115, NX116, NX117,
     NX118, NX119, NX120, NX121, NX122, NX123, NX124, NX125, NX126,
     NX127, NX128, NX129, NX130, NX131, NX132, NX133, NX134, NX135,
     NX136, NX137, NX138, NX139, NX140, NX141, NX142, NX143, NX144,
     NX145, NX146, NX147, NX148, NX149, NX150, NX151, NX152, NX153,
     NX154, NX155, NX156, NX157, NX158, NX159, NX160, NX161, NX162,
     NX163, NX164, NX165, NX166, NX167, NX168, NX169, NX170, NX171,
     NX172, NX173, NX174, NX175, NX176, NX177, NX178, NX179, NX180,
     NX181, NX182, NX183, NX184, NX185, NX186, NX187, NX188, NX189,
     NX190, NX191, NX192, NX193, NX194, NX195, NX196, NX197, NX198,
     NX199, NX200, NX201, NX202, NX203, NX204, NX205, NX206, NX207,
     NX208, NX209, NX210, NX211, NX212, NX213, NX214, NX215, NX216,
     NX217, NX218, NX219, NX220, NX221, NX222, NX223, NX224, NX225,
     NX226, NX227, NX228, NX229, NX230, NX231, NX232, NX233, NX234,
     NX235, NX236, NX237, NX238, NX239, NX240, NX241, NX242, NX243,
     NX244, NX245, NX246, NX247, NX248, NX249, NX250, NX251, NX252,
     NX253, NX254, NX255, RACK0, RACK1, RACK2, RACK3, RACK4, RACK5,
     RACK6, RACK7, RACK8, RACK9, RACK10, RACK11, RACK12, RACK13,
     RACK14, RACK15, X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, X11,
     X12, X13, X14, X15, X16, X17, X18, X19, X20, X21, X22, X23, X24,
     X25, X26, X27, X28, X29, X30, X31, X32, X33, X34, X35, X36, X37,
     X38, X39, X40, X41, X42, X43, X44, X45, X46, X47, X48, X49, X50,
     X51, X52, X53, X54, X55, X56, X57, X58, X59, X60, X61, X62, X63,
     X64, X65, X66, X67, X68, X69, X70, X71, X72, X73, X74, X75, X76,
     X77, X78, X79, X80, X81, X82, X83, X84, X85, X86, X87, X88, X89,
     X90, X91, X92, X93, X94, X95, X96, X97, X98, X99, X100, X101,
     X102, X103, X104, X105, X106, X107, X108, X109, X110, X111, X112,
     X113, X114, X115, X116, X117, X118, X119, X120, X121, X122, X123,
     X124, X125, X126, X127, X128, X129, X130, X131, X132, X133, X134,
     X135, X136, X137, X138, X139, X140, X141, X142, X143, X144, X145,
     X146, X147, X148, X149, X150, X151, X152, X153, X154, X155, X156,
     X157, X158, X159, X160, X161, X162, X163, X164, X165, X166, X167,
     X168, X169, X170, X171, X172, X173, X174, X175, X176, X177, X178,
     X179, X180, X181, X182, X183, X184, X185, X186, X187, X188, X189,
     X190, X191, X192, X193, X194, X195, X196, X197, X198, X199, X200,
     X201, X202, X203, X204, X205, X206, X207, X208, X209, X210, X211,
     X212, X213, X214, X215, X216, X217, X218, X219, X220, X221, X222,
     X223, X224, X225, X226, X227, X228, X229, X230, X231, X232, X233,
     X234, X235, X236, X237, X238, X239, X240, X241, X242, X243, X244,
     X245, X246, X247, X248, X249, X250, X251, X252, X253, X254, X255;


specify
    specparam CDS_LIBNAME  = "XB16TSMC65";
    specparam CDS_CELLNAME = "ZFBAR4";
    specparam CDS_VIEWNAME = "schematic";
endspecify

ZZFBCP I17 ( NR00, NR10, NR20, NR30, NR40, NR50, NR60, NR70, NR80,
     NR90, NR100, NR110, NR120, NR130, NR140, NR150, R00, R10, R20,
     R30, R40, R50, R60, R70, R80, R90, R100, R110, R120, R130, R140,
     R150, VDD, VSS, L00, L10, L20, L30, L40, L50, L60, L70, L80, L90,
     L100, L110, L120, L130, L140, L150, NL00, NL10, NL20, NL30, NL40,
     NL50, NL60, NL70, NL80, NL90, NL100, NL110, NL120, NL130, NL140,
     NL150, NRACK0, NRACK1, NRACK2, NRACK3, NRACK4, NRACK5, NRACK6,
     NRACK7, NRACK8, NRACK9, NRACK10, NRACK11, NRACK12, NRACK13,
     NRACK14, NRACK15, NVAL0, NX0, NX1, NX2, NX3, NX4, NX5, NX6, NX7,
     NX8, NX9, NX10, NX11, NX12, NX13, NX14, NX15, NX16, NX17, NX18,
     NX19, NX20, NX21, NX22, NX23, NX24, NX25, NX26, NX27, NX28, NX29,
     NX30, NX31, NX32, NX33, NX34, NX35, NX36, NX37, NX38, NX39, NX40,
     NX41, NX42, NX43, NX44, NX45, NX46, NX47, NX48, NX49, NX50, NX51,
     NX52, NX53, NX54, NX55, NX56, NX57, NX58, NX59, NX60, NX61, NX62,
     NX63, NX64, NX65, NX66, NX67, NX68, NX69, NX70, NX71, NX72, NX73,
     NX74, NX75, NX76, NX77, NX78, NX79, NX80, NX81, NX82, NX83, NX84,
     NX85, NX86, NX87, NX88, NX89, NX90, NX91, NX92, NX93, NX94, NX95,
     NX96, NX97, NX98, NX99, NX100, NX101, NX102, NX103, NX104, NX105,
     NX106, NX107, NX108, NX109, NX110, NX111, NX112, NX113, NX114,
     NX115, NX116, NX117, NX118, NX119, NX120, NX121, NX122, NX123,
     NX124, NX125, NX126, NX127, NX128, NX129, NX130, NX131, NX132,
     NX133, NX134, NX135, NX136, NX137, NX138, NX139, NX140, NX141,
     NX142, NX143, NX144, NX145, NX146, NX147, NX148, NX149, NX150,
     NX151, NX152, NX153, NX154, NX155, NX156, NX157, NX158, NX159,
     NX160, NX161, NX162, NX163, NX164, NX165, NX166, NX167, NX168,
     NX169, NX170, NX171, NX172, NX173, NX174, NX175, NX176, NX177,
     NX178, NX179, NX180, NX181, NX182, NX183, NX184, NX185, NX186,
     NX187, NX188, NX189, NX190, NX191, NX192, NX193, NX194, NX195,
     NX196, NX197, NX198, NX199, NX200, NX201, NX202, NX203, NX204,
     NX205, NX206, NX207, NX208, NX209, NX210, NX211, NX212, NX213,
     NX214, NX215, NX216, NX217, NX218, NX219, NX220, NX221, NX222,
     NX223, NX224, NX225, NX226, NX227, NX228, NX229, NX230, NX231,
     NX232, NX233, NX234, NX235, NX236, NX237, NX238, NX239, NX240,
     NX241, NX242, NX243, NX244, NX245, NX246, NX247, NX248, NX249,
     NX250, NX251, NX252, NX253, NX254, NX255, RACK0, RACK1, RACK2,
     RACK3, RACK4, RACK5, RACK6, RACK7, RACK8, RACK9, RACK10, RACK11,
     RACK12, RACK13, RACK14, RACK15, X0, X1, X2, X3, X4, X5, X6, X7,
     X8, X9, X10, X11, X12, X13, X14, X15, X16, X17, X18, X19, X20,
     X21, X22, X23, X24, X25, X26, X27, X28, X29, X30, X31, X32, X33,
     X34, X35, X36, X37, X38, X39, X40, X41, X42, X43, X44, X45, X46,
     X47, X48, X49, X50, X51, X52, X53, X54, X55, X56, X57, X58, X59,
     X60, X61, X62, X63, X64, X65, X66, X67, X68, X69, X70, X71, X72,
     X73, X74, X75, X76, X77, X78, X79, X80, X81, X82, X83, X84, X85,
     X86, X87, X88, X89, X90, X91, X92, X93, X94, X95, X96, X97, X98,
     X99, X100, X101, X102, X103, X104, X105, X106, X107, X108, X109,
     X110, X111, X112, X113, X114, X115, X116, X117, X118, X119, X120,
     X121, X122, X123, X124, X125, X126, X127, X128, X129, X130, X131,
     X132, X133, X134, X135, X136, X137, X138, X139, X140, X141, X142,
     X143, X144, X145, X146, X147, X148, X149, X150, X151, X152, X153,
     X154, X155, X156, X157, X158, X159, X160, X161, X162, X163, X164,
     X165, X166, X167, X168, X169, X170, X171, X172, X173, X174, X175,
     X176, X177, X178, X179, X180, X181, X182, X183, X184, X185, X186,
     X187, X188, X189, X190, X191, X192, X193, X194, X195, X196, X197,
     X198, X199, X200, X201, X202, X203, X204, X205, X206, X207, X208,
     X209, X210, X211, X212, X213, X214, X215, X216, X217, X218, X219,
     X220, X221, X222, X223, X224, X225, X226, X227, X228, X229, X230,
     X231, X232, X233, X234, X235, X236, X237, X238, X239, X240, X241,
     X242, X243, X244, X245, X246, X247, X248, X249, X250, X251, X252,
     X253, X254, X255);
ZZFBCP I20 ( NR03, NR13, NR23, NR33, NR43, NR53, NR63, NR73, NR83,
     NR93, NR103, NR113, NR123, NR133, NR143, NR153, R03, R13, R23,
     R33, R43, R53, R63, R73, R83, R93, R103, R113, R123, R133, R143,
     R153, VDD, VSS, L03, L13, L23, L33, L43, L53, L63, L73, L83, L93,
     L103, L113, L123, L133, L143, L153, NL03, NL13, NL23, NL33, NL43,
     NL53, NL63, NL73, NL83, NL93, NL103, NL113, NL123, NL133, NL143,
     NL153, NRACK0, NRACK1, NRACK2, NRACK3, NRACK4, NRACK5, NRACK6,
     NRACK7, NRACK8, NRACK9, NRACK10, NRACK11, NRACK12, NRACK13,
     NRACK14, NRACK15, NVAL3, NX0, NX1, NX2, NX3, NX4, NX5, NX6, NX7,
     NX8, NX9, NX10, NX11, NX12, NX13, NX14, NX15, NX16, NX17, NX18,
     NX19, NX20, NX21, NX22, NX23, NX24, NX25, NX26, NX27, NX28, NX29,
     NX30, NX31, NX32, NX33, NX34, NX35, NX36, NX37, NX38, NX39, NX40,
     NX41, NX42, NX43, NX44, NX45, NX46, NX47, NX48, NX49, NX50, NX51,
     NX52, NX53, NX54, NX55, NX56, NX57, NX58, NX59, NX60, NX61, NX62,
     NX63, NX64, NX65, NX66, NX67, NX68, NX69, NX70, NX71, NX72, NX73,
     NX74, NX75, NX76, NX77, NX78, NX79, NX80, NX81, NX82, NX83, NX84,
     NX85, NX86, NX87, NX88, NX89, NX90, NX91, NX92, NX93, NX94, NX95,
     NX96, NX97, NX98, NX99, NX100, NX101, NX102, NX103, NX104, NX105,
     NX106, NX107, NX108, NX109, NX110, NX111, NX112, NX113, NX114,
     NX115, NX116, NX117, NX118, NX119, NX120, NX121, NX122, NX123,
     NX124, NX125, NX126, NX127, NX128, NX129, NX130, NX131, NX132,
     NX133, NX134, NX135, NX136, NX137, NX138, NX139, NX140, NX141,
     NX142, NX143, NX144, NX145, NX146, NX147, NX148, NX149, NX150,
     NX151, NX152, NX153, NX154, NX155, NX156, NX157, NX158, NX159,
     NX160, NX161, NX162, NX163, NX164, NX165, NX166, NX167, NX168,
     NX169, NX170, NX171, NX172, NX173, NX174, NX175, NX176, NX177,
     NX178, NX179, NX180, NX181, NX182, NX183, NX184, NX185, NX186,
     NX187, NX188, NX189, NX190, NX191, NX192, NX193, NX194, NX195,
     NX196, NX197, NX198, NX199, NX200, NX201, NX202, NX203, NX204,
     NX205, NX206, NX207, NX208, NX209, NX210, NX211, NX212, NX213,
     NX214, NX215, NX216, NX217, NX218, NX219, NX220, NX221, NX222,
     NX223, NX224, NX225, NX226, NX227, NX228, NX229, NX230, NX231,
     NX232, NX233, NX234, NX235, NX236, NX237, NX238, NX239, NX240,
     NX241, NX242, NX243, NX244, NX245, NX246, NX247, NX248, NX249,
     NX250, NX251, NX252, NX253, NX254, NX255, RACK0, RACK1, RACK2,
     RACK3, RACK4, RACK5, RACK6, RACK7, RACK8, RACK9, RACK10, RACK11,
     RACK12, RACK13, RACK14, RACK15, X0, X1, X2, X3, X4, X5, X6, X7,
     X8, X9, X10, X11, X12, X13, X14, X15, X16, X17, X18, X19, X20,
     X21, X22, X23, X24, X25, X26, X27, X28, X29, X30, X31, X32, X33,
     X34, X35, X36, X37, X38, X39, X40, X41, X42, X43, X44, X45, X46,
     X47, X48, X49, X50, X51, X52, X53, X54, X55, X56, X57, X58, X59,
     X60, X61, X62, X63, X64, X65, X66, X67, X68, X69, X70, X71, X72,
     X73, X74, X75, X76, X77, X78, X79, X80, X81, X82, X83, X84, X85,
     X86, X87, X88, X89, X90, X91, X92, X93, X94, X95, X96, X97, X98,
     X99, X100, X101, X102, X103, X104, X105, X106, X107, X108, X109,
     X110, X111, X112, X113, X114, X115, X116, X117, X118, X119, X120,
     X121, X122, X123, X124, X125, X126, X127, X128, X129, X130, X131,
     X132, X133, X134, X135, X136, X137, X138, X139, X140, X141, X142,
     X143, X144, X145, X146, X147, X148, X149, X150, X151, X152, X153,
     X154, X155, X156, X157, X158, X159, X160, X161, X162, X163, X164,
     X165, X166, X167, X168, X169, X170, X171, X172, X173, X174, X175,
     X176, X177, X178, X179, X180, X181, X182, X183, X184, X185, X186,
     X187, X188, X189, X190, X191, X192, X193, X194, X195, X196, X197,
     X198, X199, X200, X201, X202, X203, X204, X205, X206, X207, X208,
     X209, X210, X211, X212, X213, X214, X215, X216, X217, X218, X219,
     X220, X221, X222, X223, X224, X225, X226, X227, X228, X229, X230,
     X231, X232, X233, X234, X235, X236, X237, X238, X239, X240, X241,
     X242, X243, X244, X245, X246, X247, X248, X249, X250, X251, X252,
     X253, X254, X255);
ZZFBCP I19 ( NR02, NR12, NR22, NR32, NR42, NR52, NR62, NR72, NR82,
     NR92, NR102, NR112, NR122, NR132, NR142, NR152, R02, R12, R22,
     R32, R42, R52, R62, R72, R82, R92, R102, R112, R122, R132, R142,
     R152, VDD, VSS, L02, L12, L22, L32, L42, L52, L62, L72, L82, L92,
     L102, L112, L122, L132, L142, L152, NL02, NL12, NL22, NL32, NL42,
     NL52, NL62, NL72, NL82, NL92, NL102, NL112, NL122, NL132, NL142,
     NL152, NRACK0, NRACK1, NRACK2, NRACK3, NRACK4, NRACK5, NRACK6,
     NRACK7, NRACK8, NRACK9, NRACK10, NRACK11, NRACK12, NRACK13,
     NRACK14, NRACK15, NVAL2, NX0, NX1, NX2, NX3, NX4, NX5, NX6, NX7,
     NX8, NX9, NX10, NX11, NX12, NX13, NX14, NX15, NX16, NX17, NX18,
     NX19, NX20, NX21, NX22, NX23, NX24, NX25, NX26, NX27, NX28, NX29,
     NX30, NX31, NX32, NX33, NX34, NX35, NX36, NX37, NX38, NX39, NX40,
     NX41, NX42, NX43, NX44, NX45, NX46, NX47, NX48, NX49, NX50, NX51,
     NX52, NX53, NX54, NX55, NX56, NX57, NX58, NX59, NX60, NX61, NX62,
     NX63, NX64, NX65, NX66, NX67, NX68, NX69, NX70, NX71, NX72, NX73,
     NX74, NX75, NX76, NX77, NX78, NX79, NX80, NX81, NX82, NX83, NX84,
     NX85, NX86, NX87, NX88, NX89, NX90, NX91, NX92, NX93, NX94, NX95,
     NX96, NX97, NX98, NX99, NX100, NX101, NX102, NX103, NX104, NX105,
     NX106, NX107, NX108, NX109, NX110, NX111, NX112, NX113, NX114,
     NX115, NX116, NX117, NX118, NX119, NX120, NX121, NX122, NX123,
     NX124, NX125, NX126, NX127, NX128, NX129, NX130, NX131, NX132,
     NX133, NX134, NX135, NX136, NX137, NX138, NX139, NX140, NX141,
     NX142, NX143, NX144, NX145, NX146, NX147, NX148, NX149, NX150,
     NX151, NX152, NX153, NX154, NX155, NX156, NX157, NX158, NX159,
     NX160, NX161, NX162, NX163, NX164, NX165, NX166, NX167, NX168,
     NX169, NX170, NX171, NX172, NX173, NX174, NX175, NX176, NX177,
     NX178, NX179, NX180, NX181, NX182, NX183, NX184, NX185, NX186,
     NX187, NX188, NX189, NX190, NX191, NX192, NX193, NX194, NX195,
     NX196, NX197, NX198, NX199, NX200, NX201, NX202, NX203, NX204,
     NX205, NX206, NX207, NX208, NX209, NX210, NX211, NX212, NX213,
     NX214, NX215, NX216, NX217, NX218, NX219, NX220, NX221, NX222,
     NX223, NX224, NX225, NX226, NX227, NX228, NX229, NX230, NX231,
     NX232, NX233, NX234, NX235, NX236, NX237, NX238, NX239, NX240,
     NX241, NX242, NX243, NX244, NX245, NX246, NX247, NX248, NX249,
     NX250, NX251, NX252, NX253, NX254, NX255, RACK0, RACK1, RACK2,
     RACK3, RACK4, RACK5, RACK6, RACK7, RACK8, RACK9, RACK10, RACK11,
     RACK12, RACK13, RACK14, RACK15, X0, X1, X2, X3, X4, X5, X6, X7,
     X8, X9, X10, X11, X12, X13, X14, X15, X16, X17, X18, X19, X20,
     X21, X22, X23, X24, X25, X26, X27, X28, X29, X30, X31, X32, X33,
     X34, X35, X36, X37, X38, X39, X40, X41, X42, X43, X44, X45, X46,
     X47, X48, X49, X50, X51, X52, X53, X54, X55, X56, X57, X58, X59,
     X60, X61, X62, X63, X64, X65, X66, X67, X68, X69, X70, X71, X72,
     X73, X74, X75, X76, X77, X78, X79, X80, X81, X82, X83, X84, X85,
     X86, X87, X88, X89, X90, X91, X92, X93, X94, X95, X96, X97, X98,
     X99, X100, X101, X102, X103, X104, X105, X106, X107, X108, X109,
     X110, X111, X112, X113, X114, X115, X116, X117, X118, X119, X120,
     X121, X122, X123, X124, X125, X126, X127, X128, X129, X130, X131,
     X132, X133, X134, X135, X136, X137, X138, X139, X140, X141, X142,
     X143, X144, X145, X146, X147, X148, X149, X150, X151, X152, X153,
     X154, X155, X156, X157, X158, X159, X160, X161, X162, X163, X164,
     X165, X166, X167, X168, X169, X170, X171, X172, X173, X174, X175,
     X176, X177, X178, X179, X180, X181, X182, X183, X184, X185, X186,
     X187, X188, X189, X190, X191, X192, X193, X194, X195, X196, X197,
     X198, X199, X200, X201, X202, X203, X204, X205, X206, X207, X208,
     X209, X210, X211, X212, X213, X214, X215, X216, X217, X218, X219,
     X220, X221, X222, X223, X224, X225, X226, X227, X228, X229, X230,
     X231, X232, X233, X234, X235, X236, X237, X238, X239, X240, X241,
     X242, X243, X244, X245, X246, X247, X248, X249, X250, X251, X252,
     X253, X254, X255);
ZZFBCP I18 ( NR01, NR11, NR21, NR31, NR41, NR51, NR61, NR71, NR81,
     NR91, NR101, NR111, NR121, NR131, NR141, NR151, R01, R11, R21,
     R31, R41, R51, R61, R71, R81, R91, R101, R111, R121, R131, R141,
     R151, VDD, VSS, L01, L11, L21, L31, L41, L51, L61, L71, L81, L91,
     L101, L111, L121, L131, L141, L151, NL01, NL11, NL21, NL31, NL41,
     NL51, NL61, NL71, NL81, NL91, NL101, NL111, NL121, NL131, NL141,
     NL151, NRACK0, NRACK1, NRACK2, NRACK3, NRACK4, NRACK5, NRACK6,
     NRACK7, NRACK8, NRACK9, NRACK10, NRACK11, NRACK12, NRACK13,
     NRACK14, NRACK15, NVAL1, NX0, NX1, NX2, NX3, NX4, NX5, NX6, NX7,
     NX8, NX9, NX10, NX11, NX12, NX13, NX14, NX15, NX16, NX17, NX18,
     NX19, NX20, NX21, NX22, NX23, NX24, NX25, NX26, NX27, NX28, NX29,
     NX30, NX31, NX32, NX33, NX34, NX35, NX36, NX37, NX38, NX39, NX40,
     NX41, NX42, NX43, NX44, NX45, NX46, NX47, NX48, NX49, NX50, NX51,
     NX52, NX53, NX54, NX55, NX56, NX57, NX58, NX59, NX60, NX61, NX62,
     NX63, NX64, NX65, NX66, NX67, NX68, NX69, NX70, NX71, NX72, NX73,
     NX74, NX75, NX76, NX77, NX78, NX79, NX80, NX81, NX82, NX83, NX84,
     NX85, NX86, NX87, NX88, NX89, NX90, NX91, NX92, NX93, NX94, NX95,
     NX96, NX97, NX98, NX99, NX100, NX101, NX102, NX103, NX104, NX105,
     NX106, NX107, NX108, NX109, NX110, NX111, NX112, NX113, NX114,
     NX115, NX116, NX117, NX118, NX119, NX120, NX121, NX122, NX123,
     NX124, NX125, NX126, NX127, NX128, NX129, NX130, NX131, NX132,
     NX133, NX134, NX135, NX136, NX137, NX138, NX139, NX140, NX141,
     NX142, NX143, NX144, NX145, NX146, NX147, NX148, NX149, NX150,
     NX151, NX152, NX153, NX154, NX155, NX156, NX157, NX158, NX159,
     NX160, NX161, NX162, NX163, NX164, NX165, NX166, NX167, NX168,
     NX169, NX170, NX171, NX172, NX173, NX174, NX175, NX176, NX177,
     NX178, NX179, NX180, NX181, NX182, NX183, NX184, NX185, NX186,
     NX187, NX188, NX189, NX190, NX191, NX192, NX193, NX194, NX195,
     NX196, NX197, NX198, NX199, NX200, NX201, NX202, NX203, NX204,
     NX205, NX206, NX207, NX208, NX209, NX210, NX211, NX212, NX213,
     NX214, NX215, NX216, NX217, NX218, NX219, NX220, NX221, NX222,
     NX223, NX224, NX225, NX226, NX227, NX228, NX229, NX230, NX231,
     NX232, NX233, NX234, NX235, NX236, NX237, NX238, NX239, NX240,
     NX241, NX242, NX243, NX244, NX245, NX246, NX247, NX248, NX249,
     NX250, NX251, NX252, NX253, NX254, NX255, RACK0, RACK1, RACK2,
     RACK3, RACK4, RACK5, RACK6, RACK7, RACK8, RACK9, RACK10, RACK11,
     RACK12, RACK13, RACK14, RACK15, X0, X1, X2, X3, X4, X5, X6, X7,
     X8, X9, X10, X11, X12, X13, X14, X15, X16, X17, X18, X19, X20,
     X21, X22, X23, X24, X25, X26, X27, X28, X29, X30, X31, X32, X33,
     X34, X35, X36, X37, X38, X39, X40, X41, X42, X43, X44, X45, X46,
     X47, X48, X49, X50, X51, X52, X53, X54, X55, X56, X57, X58, X59,
     X60, X61, X62, X63, X64, X65, X66, X67, X68, X69, X70, X71, X72,
     X73, X74, X75, X76, X77, X78, X79, X80, X81, X82, X83, X84, X85,
     X86, X87, X88, X89, X90, X91, X92, X93, X94, X95, X96, X97, X98,
     X99, X100, X101, X102, X103, X104, X105, X106, X107, X108, X109,
     X110, X111, X112, X113, X114, X115, X116, X117, X118, X119, X120,
     X121, X122, X123, X124, X125, X126, X127, X128, X129, X130, X131,
     X132, X133, X134, X135, X136, X137, X138, X139, X140, X141, X142,
     X143, X144, X145, X146, X147, X148, X149, X150, X151, X152, X153,
     X154, X155, X156, X157, X158, X159, X160, X161, X162, X163, X164,
     X165, X166, X167, X168, X169, X170, X171, X172, X173, X174, X175,
     X176, X177, X178, X179, X180, X181, X182, X183, X184, X185, X186,
     X187, X188, X189, X190, X191, X192, X193, X194, X195, X196, X197,
     X198, X199, X200, X201, X202, X203, X204, X205, X206, X207, X208,
     X209, X210, X211, X212, X213, X214, X215, X216, X217, X218, X219,
     X220, X221, X222, X223, X224, X225, X226, X227, X228, X229, X230,
     X231, X232, X233, X234, X235, X236, X237, X238, X239, X240, X241,
     X242, X243, X244, X245, X246, X247, X248, X249, X250, X251, X252,
     X253, X254, X255);

endmodule

// Library - XB16TSMC65, Cell - ZXGNAX, View - schematic
// LAST TIME SAVED: May  8 15:13:01 2023
// NETLIST TIME: May 12 11:49:59 2023
`timescale 1ns / 1ns

module ZXGNAX ( NVAE0, NVAE1, NVAE2, NVAE3, NVAE4, NVAE5, NVAE6, NVAE7,
     NVAE8, NVAE9, NVAE10, NVAE11, NVAE12, NVAE13, NVAE14, NVAE15, X0,
     X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, X11, X12, X13, X14, X15,
     X16, X17, X18, X19, X20, X21, X22, X23, X24, X25, X26, X27, X28,
     X29, X30, X31, X32, X33, X34, X35, X36, X37, X38, X39, X40, X41,
     X42, X43, X44, X45, X46, X47, X48, X49, X50, X51, X52, X53, X54,
     X55, X56, X57, X58, X59, X60, X61, X62, X63, X64, X65, X66, X67,
     X68, X69, X70, X71, X72, X73, X74, X75, X76, X77, X78, X79, X80,
     X81, X82, X83, X84, X85, X86, X87, X88, X89, X90, X91, X92, X93,
     X94, X95, X96, X97, X98, X99, X100, X101, X102, X103, X104, X105,
     X106, X107, X108, X109, X110, X111, X112, X113, X114, X115, X116,
     X117, X118, X119, X120, X121, X122, X123, X124, X125, X126, X127,
     X128, X129, X130, X131, X132, X133, X134, X135, X136, X137, X138,
     X139, X140, X141, X142, X143, X144, X145, X146, X147, X148, X149,
     X150, X151, X152, X153, X154, X155, X156, X157, X158, X159, X160,
     X161, X162, X163, X164, X165, X166, X167, X168, X169, X170, X171,
     X172, X173, X174, X175, X176, X177, X178, X179, X180, X181, X182,
     X183, X184, X185, X186, X187, X188, X189, X190, X191, X192, X193,
     X194, X195, X196, X197, X198, X199, X200, X201, X202, X203, X204,
     X205, X206, X207, X208, X209, X210, X211, X212, X213, X214, X215,
     X216, X217, X218, X219, X220, X221, X222, X223, X224, X225, X226,
     X227, X228, X229, X230, X231, X232, X233, X234, X235, X236, X237,
     X238, X239, X240, X241, X242, X243, X244, X245, X246, X247, X248,
     X249, X250, X251, X252, X253, X254, X255 );

output  NVAE0, NVAE1, NVAE2, NVAE3, NVAE4, NVAE5, NVAE6, NVAE7, NVAE8,
     NVAE9, NVAE10, NVAE11, NVAE12, NVAE13, NVAE14, NVAE15;

input  X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, X11, X12, X13, X14,
     X15, X16, X17, X18, X19, X20, X21, X22, X23, X24, X25, X26, X27,
     X28, X29, X30, X31, X32, X33, X34, X35, X36, X37, X38, X39, X40,
     X41, X42, X43, X44, X45, X46, X47, X48, X49, X50, X51, X52, X53,
     X54, X55, X56, X57, X58, X59, X60, X61, X62, X63, X64, X65, X66,
     X67, X68, X69, X70, X71, X72, X73, X74, X75, X76, X77, X78, X79,
     X80, X81, X82, X83, X84, X85, X86, X87, X88, X89, X90, X91, X92,
     X93, X94, X95, X96, X97, X98, X99, X100, X101, X102, X103, X104,
     X105, X106, X107, X108, X109, X110, X111, X112, X113, X114, X115,
     X116, X117, X118, X119, X120, X121, X122, X123, X124, X125, X126,
     X127, X128, X129, X130, X131, X132, X133, X134, X135, X136, X137,
     X138, X139, X140, X141, X142, X143, X144, X145, X146, X147, X148,
     X149, X150, X151, X152, X153, X154, X155, X156, X157, X158, X159,
     X160, X161, X162, X163, X164, X165, X166, X167, X168, X169, X170,
     X171, X172, X173, X174, X175, X176, X177, X178, X179, X180, X181,
     X182, X183, X184, X185, X186, X187, X188, X189, X190, X191, X192,
     X193, X194, X195, X196, X197, X198, X199, X200, X201, X202, X203,
     X204, X205, X206, X207, X208, X209, X210, X211, X212, X213, X214,
     X215, X216, X217, X218, X219, X220, X221, X222, X223, X224, X225,
     X226, X227, X228, X229, X230, X231, X232, X233, X234, X235, X236,
     X237, X238, X239, X240, X241, X242, X243, X244, X245, X246, X247,
     X248, X249, X250, X251, X252, X253, X254, X255;


specify
    specparam CDS_LIBNAME  = "XB16TSMC65";
    specparam CDS_CELLNAME = "ZXGNAX";
    specparam CDS_VIEWNAME = "schematic";
endspecify

INVXB1 I176 ( NVAE15, cds_globals.vdd_, cds_globals.gnd_, net0213);
INVXB1 I175 ( net0213, cds_globals.vdd_, cds_globals.gnd_, net0211);
INVXB1 I174 ( NVAE14, cds_globals.vdd_, cds_globals.gnd_, net0191);
INVXB1 I173 ( net0191, cds_globals.vdd_, cds_globals.gnd_, net0230);
INVXB1 I172 ( NVAE13, cds_globals.vdd_, cds_globals.gnd_, net0193);
INVXB1 I171 ( net0193, cds_globals.vdd_, cds_globals.gnd_, net0233);
INVXB1 I170 ( NVAE12, cds_globals.vdd_, cds_globals.gnd_, net0179);
INVXB1 I169 ( net0179, cds_globals.vdd_, cds_globals.gnd_, net0195);
INVXB1 I168 ( NVAE11, cds_globals.vdd_, cds_globals.gnd_, net0210);
INVXB1 I167 ( net0210, cds_globals.vdd_, cds_globals.gnd_, net0203);
INVXB1 I166 ( NVAE10, cds_globals.vdd_, cds_globals.gnd_, net0223);
INVXB1 I165 ( net0223, cds_globals.vdd_, cds_globals.gnd_, net0232);
INVXB1 I164 ( NVAE9, cds_globals.vdd_, cds_globals.gnd_, net0206);
INVXB1 I163 ( net0206, cds_globals.vdd_, cds_globals.gnd_, net0231);
INVXB1 I162 ( NVAE8, cds_globals.vdd_, cds_globals.gnd_, net0192);
INVXB1 I161 ( net0192, cds_globals.vdd_, cds_globals.gnd_, net0228);
INVXB1 I160 ( NVAE7, cds_globals.vdd_, cds_globals.gnd_, net0189);
INVXB1 I159 ( net0189, cds_globals.vdd_, cds_globals.gnd_, net0161);
INVXB1 I158 ( NVAE6, cds_globals.vdd_, cds_globals.gnd_, net0177);
INVXB1 I157 ( net0177, cds_globals.vdd_, cds_globals.gnd_, net0181);
INVXB1 I156 ( NVAE5, cds_globals.vdd_, cds_globals.gnd_, net0215);
INVXB1 I155 ( net0215, cds_globals.vdd_, cds_globals.gnd_, net0209);
INVXB1 I154 ( NVAE4, cds_globals.vdd_, cds_globals.gnd_, net0175);
INVXB1 I153 ( net0175, cds_globals.vdd_, cds_globals.gnd_, net0222);
INVXB1 I152 ( NVAE3, cds_globals.vdd_, cds_globals.gnd_, net0212);
INVXB1 I151 ( net0212, cds_globals.vdd_, cds_globals.gnd_, net0229);
INVXB1 I150 ( NVAE2, cds_globals.vdd_, cds_globals.gnd_, net0188);
INVXB1 I149 ( net0188, cds_globals.vdd_, cds_globals.gnd_, net0220);
INVXB1 I148 ( NVAE1, cds_globals.vdd_, cds_globals.gnd_, net093);
INVXB1 I147 ( net093, cds_globals.vdd_, cds_globals.gnd_, net094);
INVXB1 I146 ( NVAE0, cds_globals.vdd_, cds_globals.gnd_, net095);
INVXB1 I145 ( net095, cds_globals.vdd_, cds_globals.gnd_, net0156);
INVXB1 I144 ( net0151, cds_globals.vdd_, cds_globals.gnd_, net0160);
INVXB1 I143 ( net0166, cds_globals.vdd_, cds_globals.gnd_, net0158);
INVXB1 I142 ( net0169, cds_globals.vdd_, cds_globals.gnd_, net0145);
INVXB1 I141 ( net0143, cds_globals.vdd_, cds_globals.gnd_, net0173);
INVXB1 I135 ( net036, cds_globals.vdd_, cds_globals.gnd_, net069);
INVXB1 I134 ( net0144, cds_globals.vdd_, cds_globals.gnd_, net070);
INVXB1 I133 ( net0154, cds_globals.vdd_, cds_globals.gnd_, net071);
INVXB1 I132 ( net035, cds_globals.vdd_, cds_globals.gnd_, net072);
INVXB1 I126 ( net0168, cds_globals.vdd_, cds_globals.gnd_, net073);
INVXB1 I125 ( net0174, cds_globals.vdd_, cds_globals.gnd_, net074);
INVXB1 I124 ( net0134, cds_globals.vdd_, cds_globals.gnd_, net075);
INVXB1 I123 ( net0172, cds_globals.vdd_, cds_globals.gnd_, net076);
INVXB1 I117 ( net0146, cds_globals.vdd_, cds_globals.gnd_, net077);
INVXB1 I116 ( net0133, cds_globals.vdd_, cds_globals.gnd_, net078);
INVXB1 I115 ( net0157, cds_globals.vdd_, cds_globals.gnd_, net079);
INVXB1 I114 ( net0171, cds_globals.vdd_, cds_globals.gnd_, net080);
INVXB1 I108 ( net0140, cds_globals.vdd_, cds_globals.gnd_, net081);
INVXB1 I107 ( net0148, cds_globals.vdd_, cds_globals.gnd_, net082);
INVXB1 I106 ( net0137, cds_globals.vdd_, cds_globals.gnd_, net083);
INVXB1 I105 ( net0152, cds_globals.vdd_, cds_globals.gnd_, net084);
INVXB1 I99 ( net0138, cds_globals.vdd_, cds_globals.gnd_, net085);
INVXB1 I98 ( net0167, cds_globals.vdd_, cds_globals.gnd_, net086);
INVXB1 I97 ( net0170, cds_globals.vdd_, cds_globals.gnd_, net087);
INVXB1 I96 ( net0132, cds_globals.vdd_, cds_globals.gnd_, net088);
INVXB1 I90 ( net0164, cds_globals.vdd_, cds_globals.gnd_, net089);
INVXB1 I89 ( net0142, cds_globals.vdd_, cds_globals.gnd_, net090);
INVXB1 I88 ( net0159, cds_globals.vdd_, cds_globals.gnd_, net091);
INVXB1 I87 ( net0129, cds_globals.vdd_, cds_globals.gnd_, net092);
INVXB1 I81 ( net020, cds_globals.vdd_, cds_globals.gnd_, net037);
INVXB1 I80 ( net02, cds_globals.vdd_, cds_globals.gnd_, net038);
INVXB1 I79 ( net01, cds_globals.vdd_, cds_globals.gnd_, net039);
INVXB1 I78 ( net019, cds_globals.vdd_, cds_globals.gnd_, net040);
INVXB1 I72 ( net022, cds_globals.vdd_, cds_globals.gnd_, net041);
INVXB1 I71 ( net04, cds_globals.vdd_, cds_globals.gnd_, net042);
INVXB1 I70 ( net03, cds_globals.vdd_, cds_globals.gnd_, net043);
INVXB1 I68 ( net021, cds_globals.vdd_, cds_globals.gnd_, net044);
INVXB1 I59 ( net024, cds_globals.vdd_, cds_globals.gnd_, net045);
INVXB1 I58 ( net06, cds_globals.vdd_, cds_globals.gnd_, net046);
INVXB1 I57 ( net05, cds_globals.vdd_, cds_globals.gnd_, net047);
INVXB1 I56 ( net023, cds_globals.vdd_, cds_globals.gnd_, net048);
INVXB1 I50 ( net026, cds_globals.vdd_, cds_globals.gnd_, net049);
INVXB1 I49 ( net08, cds_globals.vdd_, cds_globals.gnd_, net050);
INVXB1 I48 ( net07, cds_globals.vdd_, cds_globals.gnd_, net051);
INVXB1 I47 ( net025, cds_globals.vdd_, cds_globals.gnd_, net052);
INVXB1 I41 ( net028, cds_globals.vdd_, cds_globals.gnd_, net053);
INVXB1 I40 ( net010, cds_globals.vdd_, cds_globals.gnd_, net054);
INVXB1 I39 ( net09, cds_globals.vdd_, cds_globals.gnd_, net055);
INVXB1 I38 ( net027, cds_globals.vdd_, cds_globals.gnd_, net056);
INVXB1 I32 ( net030, cds_globals.vdd_, cds_globals.gnd_, net057);
INVXB1 I31 ( net012, cds_globals.vdd_, cds_globals.gnd_, net058);
INVXB1 I30 ( net011, cds_globals.vdd_, cds_globals.gnd_, net059);
INVXB1 I29 ( net029, cds_globals.vdd_, cds_globals.gnd_, net060);
INVXB1 I12 ( net015, cds_globals.vdd_, cds_globals.gnd_, net067);
INVXB1 I62 ( net1, cds_globals.vdd_, cds_globals.gnd_, net2);
INVXB1 I23 ( net032, cds_globals.vdd_, cds_globals.gnd_, net061);
INVXB1 I22 ( net014, cds_globals.vdd_, cds_globals.gnd_, net062);
INVXB1 I21 ( net013, cds_globals.vdd_, cds_globals.gnd_, net063);
INVXB1 I65 ( net6, cds_globals.vdd_, cds_globals.gnd_, net7);
INVXB1 I20 ( net031, cds_globals.vdd_, cds_globals.gnd_, net064);
INVXB1 I66 ( net5, cds_globals.vdd_, cds_globals.gnd_, net8);
INVXB1 I69 ( net4, cds_globals.vdd_, cds_globals.gnd_, net9);
INVXB1 I14 ( net034, cds_globals.vdd_, cds_globals.gnd_, net065);
INVXB1 I13 ( net016, cds_globals.vdd_, cds_globals.gnd_, net066);
INVXB1 I11 ( net033, cds_globals.vdd_, cds_globals.gnd_, net068);
NR4XB1 I140 ( net0158, cds_globals.vdd_, cds_globals.gnd_, X79, X95,
     X111, X127);
NR4XB1 I139 ( net0145, cds_globals.vdd_, cds_globals.gnd_, X143, X159,
     X175, X191);
NR4XB1 I138 ( net0173, cds_globals.vdd_, cds_globals.gnd_, X207, X223,
     X239, X255);
NR4XB1 I137 ( net0160, cds_globals.vdd_, cds_globals.gnd_, X15, X31,
     X47, X63);
NR4XB1 I136 ( net0211, cds_globals.vdd_, cds_globals.gnd_, net0151,
     net0166, net0169, net0143);
NR4XB1 I131 ( net070, cds_globals.vdd_, cds_globals.gnd_, X78, X94,
     X110, X126);
NR4XB1 I130 ( net071, cds_globals.vdd_, cds_globals.gnd_, X142, X158,
     X174, X190);
NR4XB1 I129 ( net072, cds_globals.vdd_, cds_globals.gnd_, X206, X222,
     X238, X254);
NR4XB1 I128 ( net069, cds_globals.vdd_, cds_globals.gnd_, X14, X30,
     X46, X62);
NR4XB1 I127 ( net0230, cds_globals.vdd_, cds_globals.gnd_, net036,
     net0144, net0154, net035);
NR4XB1 I122 ( net074, cds_globals.vdd_, cds_globals.gnd_, X77, X93,
     X109, X125);
NR4XB1 I121 ( net075, cds_globals.vdd_, cds_globals.gnd_, X141, X157,
     X173, X189);
NR4XB1 I120 ( net076, cds_globals.vdd_, cds_globals.gnd_, X205, X221,
     X237, X253);
NR4XB1 I119 ( net073, cds_globals.vdd_, cds_globals.gnd_, X13, X29,
     X45, X61);
NR4XB1 I118 ( net0233, cds_globals.vdd_, cds_globals.gnd_, net0168,
     net0174, net0134, net0172);
NR4XB1 I113 ( net078, cds_globals.vdd_, cds_globals.gnd_, X76, X92,
     X108, X124);
NR4XB1 I112 ( net079, cds_globals.vdd_, cds_globals.gnd_, X140, X156,
     X172, X188);
NR4XB1 I111 ( net080, cds_globals.vdd_, cds_globals.gnd_, X204, X220,
     X236, X252);
NR4XB1 I110 ( net077, cds_globals.vdd_, cds_globals.gnd_, X12, X28,
     X44, X60);
NR4XB1 I109 ( net0195, cds_globals.vdd_, cds_globals.gnd_, net0146,
     net0133, net0157, net0171);
NR4XB1 I104 ( net082, cds_globals.vdd_, cds_globals.gnd_, X75, X91,
     X107, X123);
NR4XB1 I103 ( net083, cds_globals.vdd_, cds_globals.gnd_, X139, X155,
     X171, X187);
NR4XB1 I102 ( net084, cds_globals.vdd_, cds_globals.gnd_, X203, X219,
     X235, X251);
NR4XB1 I101 ( net081, cds_globals.vdd_, cds_globals.gnd_, X11, X27,
     X43, X59);
NR4XB1 I100 ( net0203, cds_globals.vdd_, cds_globals.gnd_, net0140,
     net0148, net0137, net0152);
NR4XB1 I95 ( net086, cds_globals.vdd_, cds_globals.gnd_, X74, X90,
     X106, X122);
NR4XB1 I94 ( net087, cds_globals.vdd_, cds_globals.gnd_, X138, X154,
     X170, X186);
NR4XB1 I93 ( net088, cds_globals.vdd_, cds_globals.gnd_, X202, X218,
     X234, X250);
NR4XB1 I92 ( net085, cds_globals.vdd_, cds_globals.gnd_, X10, X26, X42,
     X58);
NR4XB1 I91 ( net0232, cds_globals.vdd_, cds_globals.gnd_, net0138,
     net0167, net0170, net0132);
NR4XB1 I86 ( net090, cds_globals.vdd_, cds_globals.gnd_, X73, X89,
     X105, X121);
NR4XB1 I85 ( net091, cds_globals.vdd_, cds_globals.gnd_, X137, X153,
     X169, X185);
NR4XB1 I84 ( net092, cds_globals.vdd_, cds_globals.gnd_, X201, X217,
     X233, X249);
NR4XB1 I83 ( net089, cds_globals.vdd_, cds_globals.gnd_, X9, X25, X41,
     X57);
NR4XB1 I82 ( net0231, cds_globals.vdd_, cds_globals.gnd_, net0164,
     net0142, net0159, net0129);
NR4XB1 I77 ( net038, cds_globals.vdd_, cds_globals.gnd_, X72, X88,
     X104, X120);
NR4XB1 I76 ( net039, cds_globals.vdd_, cds_globals.gnd_, X136, X152,
     X168, X184);
NR4XB1 I75 ( net040, cds_globals.vdd_, cds_globals.gnd_, X200, X216,
     X232, X248);
NR4XB1 I74 ( net037, cds_globals.vdd_, cds_globals.gnd_, X8, X24, X40,
     X56);
NR4XB1 I73 ( net0228, cds_globals.vdd_, cds_globals.gnd_, net020,
     net02, net01, net019);
NR4XB1 I67 ( net042, cds_globals.vdd_, cds_globals.gnd_, X71, X87,
     X103, X119);
NR4XB1 I64 ( net043, cds_globals.vdd_, cds_globals.gnd_, X135, X151,
     X167, X183);
NR4XB1 I63 ( net044, cds_globals.vdd_, cds_globals.gnd_, X199, X215,
     X231, X247);
NR4XB1 I61 ( net041, cds_globals.vdd_, cds_globals.gnd_, X7, X23, X39,
     X55);
NR4XB1 I60 ( net0161, cds_globals.vdd_, cds_globals.gnd_, net022,
     net04, net03, net021);
NR4XB1 I55 ( net046, cds_globals.vdd_, cds_globals.gnd_, X70, X86,
     X102, X118);
NR4XB1 I54 ( net047, cds_globals.vdd_, cds_globals.gnd_, X134, X150,
     X166, X182);
NR4XB1 I53 ( net048, cds_globals.vdd_, cds_globals.gnd_, X198, X214,
     X230, X246);
NR4XB1 I52 ( net045, cds_globals.vdd_, cds_globals.gnd_, X6, X22, X38,
     X54);
NR4XB1 I51 ( net0181, cds_globals.vdd_, cds_globals.gnd_, net024,
     net06, net05, net023);
NR4XB1 I46 ( net050, cds_globals.vdd_, cds_globals.gnd_, X69, X85,
     X101, X117);
NR4XB1 I45 ( net051, cds_globals.vdd_, cds_globals.gnd_, X133, X149,
     X165, X181);
NR4XB1 I44 ( net052, cds_globals.vdd_, cds_globals.gnd_, X197, X213,
     X229, X245);
NR4XB1 I43 ( net049, cds_globals.vdd_, cds_globals.gnd_, X5, X21, X37,
     X53);
NR4XB1 I42 ( net0209, cds_globals.vdd_, cds_globals.gnd_, net026,
     net08, net07, net025);
NR4XB1 I37 ( net054, cds_globals.vdd_, cds_globals.gnd_, X68, X84,
     X100, X116);
NR4XB1 I36 ( net055, cds_globals.vdd_, cds_globals.gnd_, X132, X148,
     X164, X180);
NR4XB1 I35 ( net056, cds_globals.vdd_, cds_globals.gnd_, X196, X212,
     X228, X244);
NR4XB1 I34 ( net053, cds_globals.vdd_, cds_globals.gnd_, X4, X20, X36,
     X52);
NR4XB1 I33 ( net0222, cds_globals.vdd_, cds_globals.gnd_, net028,
     net010, net09, net027);
NR4XB1 I28 ( net058, cds_globals.vdd_, cds_globals.gnd_, X67, X83, X99,
     X115);
NR4XB1 I27 ( net059, cds_globals.vdd_, cds_globals.gnd_, X131, X147,
     X163, X179);
NR4XB1 I26 ( net060, cds_globals.vdd_, cds_globals.gnd_, X195, X211,
     X227, X243);
NR4XB1 I25 ( net057, cds_globals.vdd_, cds_globals.gnd_, X3, X19, X35,
     X51);
NR4XB1 I24 ( net0229, cds_globals.vdd_, cds_globals.gnd_, net030,
     net012, net011, net029);
NR4XB1 I8 ( net068, cds_globals.vdd_, cds_globals.gnd_, X193, X209,
     X225, X241);
NR4XB1 I9 ( net067, cds_globals.vdd_, cds_globals.gnd_, X129, X145,
     X161, X177);
NR4XB1 I7 ( net065, cds_globals.vdd_, cds_globals.gnd_, X1, X17, X33,
     X49);
NR4XB1 I3 ( net9, cds_globals.vdd_, cds_globals.gnd_, X192, X208, X224,
     X240);
NR4XB1 I19 ( net062, cds_globals.vdd_, cds_globals.gnd_, X66, X82, X98,
     X114);
NR4XB1 I6 ( net094, cds_globals.vdd_, cds_globals.gnd_, net034, net016,
     net015, net033);
NR4XB1 I18 ( net063, cds_globals.vdd_, cds_globals.gnd_, X130, X146,
     X162, X178);
NR4XB1 I2 ( net8, cds_globals.vdd_, cds_globals.gnd_, X128, X144, X160,
     X176);
NR4XB1 I17 ( net064, cds_globals.vdd_, cds_globals.gnd_, X194, X210,
     X226, X242);
NR4XB1 I5 ( net0156, cds_globals.vdd_, cds_globals.gnd_, net1, net6,
     net5, net4);
NR4XB1 I16 ( net061, cds_globals.vdd_, cds_globals.gnd_, X2, X18, X34,
     X50);
NR4XB1 I15 ( net0220, cds_globals.vdd_, cds_globals.gnd_, net032,
     net014, net013, net031);
NR4XB1 I1 ( net7, cds_globals.vdd_, cds_globals.gnd_, X64, X80, X96,
     X112);
NR4XB1 I0 ( net2, cds_globals.vdd_, cds_globals.gnd_, X0, X16, X32,
     X48);
NR4XB1 I10 ( net066, cds_globals.vdd_, cds_globals.gnd_, X65, X81, X97,
     X113);

endmodule

// Library - XB16TSMC65, Cell - ZLCKAO, View - schematic
// LAST TIME SAVED: May  8 15:13:02 2023
// NETLIST TIME: May 12 11:49:59 2023
`timescale 1ns / 1ns

module ZLCKAO ( NLACK0, NLACK1, NLACK2, NLACK3, NLACK4, NLACK5, NLACK6,
     NLACK7, NLACK8, NLACK9, NLACK10, NLACK11, NLACK12, NLACK13,
     NLACK14, NLACK15, NS0, NS1, NS2, NS3, NS4, NS5, NS6, NS7, NS8,
     NS9, NS10, NS11, NS12, NS13, NS14, NS15, Rval );

output  NLACK0, NLACK1, NLACK2, NLACK3, NLACK4, NLACK5, NLACK6, NLACK7,
     NLACK8, NLACK9, NLACK10, NLACK11, NLACK12, NLACK13, NLACK14,
     NLACK15;

input  NS0, NS1, NS2, NS3, NS4, NS5, NS6, NS7, NS8, NS9, NS10, NS11,
     NS12, NS13, NS14, NS15, Rval;


specify
    specparam CDS_LIBNAME  = "XB16TSMC65";
    specparam CDS_CELLNAME = "ZLCKAO";
    specparam CDS_VIEWNAME = "schematic";
endspecify

CEL2XB1 I269 ( NLACK0, cds_globals.vdd_, cds_globals.gnd_, NS0, Rval);
CEL2XB1 I279 ( NLACK15, cds_globals.vdd_, cds_globals.gnd_, NS15,
     Rval);
CEL2XB1 I278 ( NLACK5, cds_globals.vdd_, cds_globals.gnd_, NS5, Rval);
CEL2XB1 I280 ( NLACK14, cds_globals.vdd_, cds_globals.gnd_, NS14,
     Rval);
CEL2XB1 I271 ( NLACK2, cds_globals.vdd_, cds_globals.gnd_, NS2, Rval);
CEL2XB1 I270 ( NLACK1, cds_globals.vdd_, cds_globals.gnd_, NS1, Rval);
CEL2XB1 I275 ( NLACK8, cds_globals.vdd_, cds_globals.gnd_, NS8, Rval);
CEL2XB1 I274 ( NLACK9, cds_globals.vdd_, cds_globals.gnd_, NS9, Rval);
CEL2XB1 I283 ( NLACK11, cds_globals.vdd_, cds_globals.gnd_, NS11,
     Rval);
CEL2XB1 I282 ( NLACK12, cds_globals.vdd_, cds_globals.gnd_, NS12,
     Rval);
CEL2XB1 I281 ( NLACK13, cds_globals.vdd_, cds_globals.gnd_, NS13,
     Rval);
CEL2XB1 I277 ( NLACK6, cds_globals.vdd_, cds_globals.gnd_, NS6, Rval);
CEL2XB1 I276 ( NLACK7, cds_globals.vdd_, cds_globals.gnd_, NS7, Rval);
CEL2XB1 I273 ( NLACK4, cds_globals.vdd_, cds_globals.gnd_, NS4, Rval);
CEL2XB1 I272 ( NLACK3, cds_globals.vdd_, cds_globals.gnd_, NS3, Rval);
CEL2XB1 I284 ( NLACK10, cds_globals.vdd_, cds_globals.gnd_, NS10,
     Rval);

endmodule


// Library - XB16TSMC65, Cell - ZCLAR4, View - schematic
// LAST TIME SAVED: May  8 15:13:02 2023
// NETLIST TIME: May 12 11:49:59 2023
`timescale 1ns / 1ns

module ZCLAR4 ( NR00, NR01, NR02, NR03, NR10, NR11, NR12, NR13, NR20,
     NR21, NR22, NR23, NR30, NR31, NR32, NR33, NR40, NR41, NR42, NR43,
     NR50, NR51, NR52, NR53, NR60, NR61, NR62, NR63, NR70, NR71, NR72,
     NR73, NR80, NR81, NR82, NR83, NR90, NR91, NR92, NR93, NR100,
     NR101, NR102, NR103, NR110, NR111, NR112, NR113, NR120, NR121,
     NR122, NR123, NR130, NR131, NR132, NR133, NR140, NR141, NR142,
     NR143, NR150, NR151, NR152, NR153, R00, R01, R02, R03, R10, R11,
     R12, R13, R20, R21, R22, R23, R30, R31, R32, R33, R40, R41, R42,
     R43, R50, R51, R52, R53, R60, R61, R62, R63, R70, R71, R72, R73,
     R80, R81, R82, R83, R90, R91, R92, R93, R100, R101, R102, R103,
     R110, R111, R112, R113, R120, R121, R122, R123, R130, R131, R132,
     R133, R140, R141, R142, R143, R150, R151, R152, R153, VDD, VSS,
     NVAL0, NVAL1, NVAL2, NVAL3, RACK0, RACK1, RACK2, RACK3, RACK4,
     RACK5, RACK6, RACK7, RACK8, RACK9, RACK10, RACK11, RACK12, RACK13,
     RACK14, RACK15 );

inout  NR00, NR01, NR02, NR03, NR10, NR11, NR12, NR13, NR20, NR21,
     NR22, NR23, NR30, NR31, NR32, NR33, NR40, NR41, NR42, NR43, NR50,
     NR51, NR52, NR53, NR60, NR61, NR62, NR63, NR70, NR71, NR72, NR73,
     NR80, NR81, NR82, NR83, NR90, NR91, NR92, NR93, NR100, NR101,
     NR102, NR103, NR110, NR111, NR112, NR113, NR120, NR121, NR122,
     NR123, NR130, NR131, NR132, NR133, NR140, NR141, NR142, NR143,
     NR150, NR151, NR152, NR153, R00, R01, R02, R03, R10, R11, R12,
     R13, R20, R21, R22, R23, R30, R31, R32, R33, R40, R41, R42, R43,
     R50, R51, R52, R53, R60, R61, R62, R63, R70, R71, R72, R73, R80,
     R81, R82, R83, R90, R91, R92, R93, R100, R101, R102, R103, R110,
     R111, R112, R113, R120, R121, R122, R123, R130, R131, R132, R133,
     R140, R141, R142, R143, R150, R151, R152, R153, VDD, VSS;

input  NVAL0, NVAL1, NVAL2, NVAL3, RACK0, RACK1, RACK2, RACK3, RACK4,
     RACK5, RACK6, RACK7, RACK8, RACK9, RACK10, RACK11, RACK12, RACK13,
     RACK14, RACK15;


specify
    specparam CDS_LIBNAME  = "XB16TSMC65";
    specparam CDS_CELLNAME = "ZCLAR4";
    specparam CDS_VIEWNAME = "schematic";
endspecify

CLSAXB1 I31 ( NR150, NR151, R150, R151, VDD, VSS, NVAL0, NVAL1,
     RACK15);
CLSAXB1 I30 ( NR152, NR153, R152, R153, VDD, VSS, NVAL2, NVAL3,
     RACK15);
CLSAXB1 I29 ( NR102, NR103, R102, R103, VDD, VSS, NVAL2, NVAL3,
     RACK10);
CLSAXB1 I28 ( NR100, NR101, R100, R101, VDD, VSS, NVAL0, NVAL1,
     RACK10);
CLSAXB1 I27 ( NR110, NR111, R110, R111, VDD, VSS, NVAL0, NVAL1,
     RACK11);
CLSAXB1 I26 ( NR112, NR113, R112, R113, VDD, VSS, NVAL2, NVAL3,
     RACK11);
CLSAXB1 I25 ( NR120, NR121, R120, R121, VDD, VSS, NVAL0, NVAL1,
     RACK12);
CLSAXB1 I24 ( NR122, NR123, R122, R123, VDD, VSS, NVAL2, NVAL3,
     RACK12);
CLSAXB1 I23 ( NR130, NR131, R130, R131, VDD, VSS, NVAL0, NVAL1,
     RACK13);
CLSAXB1 I22 ( NR132, NR133, R132, R133, VDD, VSS, NVAL2, NVAL3,
     RACK13);
CLSAXB1 I21 ( NR140, NR141, R140, R141, VDD, VSS, NVAL0, NVAL1,
     RACK14);
CLSAXB1 I20 ( NR142, NR143, R142, R143, VDD, VSS, NVAL2, NVAL3,
     RACK14);
CLSAXB1 I19 ( NR52, NR53, R52, R53, VDD, VSS, NVAL2, NVAL3, RACK5);
CLSAXB1 I18 ( NR50, NR51, R50, R51, VDD, VSS, NVAL0, NVAL1, RACK5);
CLSAXB1 I17 ( NR60, NR61, R60, R61, VDD, VSS, NVAL0, NVAL1, RACK6);
CLSAXB1 I16 ( NR62, NR63, R62, R63, VDD, VSS, NVAL2, NVAL3, RACK6);
CLSAXB1 I15 ( NR70, NR71, R70, R71, VDD, VSS, NVAL0, NVAL1, RACK7);
CLSAXB1 I14 ( NR72, NR73, R72, R73, VDD, VSS, NVAL2, NVAL3, RACK7);
CLSAXB1 I13 ( NR80, NR81, R80, R81, VDD, VSS, NVAL0, NVAL1, RACK8);
CLSAXB1 I12 ( NR82, NR83, R82, R83, VDD, VSS, NVAL2, NVAL3, RACK8);
CLSAXB1 I11 ( NR90, NR91, R90, R91, VDD, VSS, NVAL0, NVAL1, RACK9);
CLSAXB1 I10 ( NR92, NR93, R92, R93, VDD, VSS, NVAL2, NVAL3, RACK9);
CLSAXB1 I9 ( NR40, NR41, R40, R41, VDD, VSS, NVAL0, NVAL1, RACK4);
CLSAXB1 I8 ( NR42, NR43, R42, R43, VDD, VSS, NVAL2, NVAL3, RACK4);
CLSAXB1 I7 ( NR20, NR21, R20, R21, VDD, VSS, NVAL0, NVAL1, RACK2);
CLSAXB1 I6 ( NR30, NR31, R30, R31, VDD, VSS, NVAL0, NVAL1, RACK3);
CLSAXB1 I5 ( NR32, NR33, R32, R33, VDD, VSS, NVAL2, NVAL3, RACK3);
CLSAXB1 I4 ( NR22, NR23, R22, R23, VDD, VSS, NVAL2, NVAL3, RACK2);
CLSAXB1 I3 ( NR10, NR11, R10, R11, VDD, VSS, NVAL0, NVAL1, RACK1);
CLSAXB1 I2 ( NR12, NR13, R12, R13, VDD, VSS, NVAL2, NVAL3, RACK1);
CLSAXB1 I1 ( NR02, NR03, R02, R03, VDD, VSS, NVAL2, NVAL3, RACK0);
CLSAXB1 I0 ( NR00, NR01, R00, R01, VDD, VSS, NVAL0, NVAL1, RACK0);

endmodule





// Library - XB16TSMC65, Cell - ZRVLAR, View - schematic
// LAST TIME SAVED: May  8 15:13:02 2023
// NETLIST TIME: May 12 11:49:58 2023
`timescale 1ns / 1ns

module ZRVLAR ( Rval, nRd00, nRd01, nRd02, nRd03, nRd10, nRd11, nRd12,
     nRd13, nRd20, nRd21, nRd22, nRd23, nRd30, nRd31, nRd32, nRd33,
     nRd40, nRd41, nRd42, nRd43, nRd50, nRd51, nRd52, nRd53, nRd60,
     nRd61, nRd62, nRd63, nRd70, nRd71, nRd72, nRd73, nRd80, nRd81,
     nRd82, nRd83, nRd90, nRd91, nRd92, nRd93, nRd100, nRd101, nRd102,
     nRd103, nRd110, nRd111, nRd112, nRd113, nRd120, nRd121, nRd122,
     nRd123, nRd130, nRd131, nRd132, nRd133, nRd140, nRd141, nRd142,
     nRd143, nRd150, nRd151, nRd152, nRd153 );

output  Rval;

input  nRd00, nRd01, nRd02, nRd03, nRd10, nRd11, nRd12, nRd13, nRd20,
     nRd21, nRd22, nRd23, nRd30, nRd31, nRd32, nRd33, nRd40, nRd41,
     nRd42, nRd43, nRd50, nRd51, nRd52, nRd53, nRd60, nRd61, nRd62,
     nRd63, nRd70, nRd71, nRd72, nRd73, nRd80, nRd81, nRd82, nRd83,
     nRd90, nRd91, nRd92, nRd93, nRd100, nRd101, nRd102, nRd103,
     nRd110, nRd111, nRd112, nRd113, nRd120, nRd121, nRd122, nRd123,
     nRd130, nRd131, nRd132, nRd133, nRd140, nRd141, nRd142, nRd143,
     nRd150, nRd151, nRd152, nRd153;


specify
    specparam CDS_LIBNAME  = "XB16TSMC65";
    specparam CDS_CELLNAME = "ZRVLAR";
    specparam CDS_VIEWNAME = "schematic";
endspecify

NR4XB1 I242 ( net027, cds_globals.vdd_, cds_globals.gnd_, net037,
     net012, net011, net028);
NR4XB1 I238 ( net029, cds_globals.vdd_, cds_globals.gnd_, nRd123,
     nRd133, nRd143, nRd153);
NR4XB1 I236 ( net032, cds_globals.vdd_, cds_globals.gnd_, nRd83, nRd93,
     nRd103, nRd113);
NR4XB1 I230 ( net035, cds_globals.vdd_, cds_globals.gnd_, nRd43, nRd53,
     nRd63, nRd73);
NR4XB1 I228 ( net038, cds_globals.vdd_, cds_globals.gnd_, nRd03, nRd13,
     nRd23, nRd33);
NR4XB1 I224 ( net040, cds_globals.vdd_, cds_globals.gnd_, net022,
     net047, net013, net041);
NR4XB1 I220 ( net042, cds_globals.vdd_, cds_globals.gnd_, nRd122,
     nRd132, nRd142, nRd152);
NR4XB1 I218 ( net045, cds_globals.vdd_, cds_globals.gnd_, nRd82, nRd92,
     nRd102, nRd112);
NR4XB1 I212 ( net048, cds_globals.vdd_, cds_globals.gnd_, nRd42, nRd52,
     nRd62, nRd72);
NR4XB1 I210 ( net051, cds_globals.vdd_, cds_globals.gnd_, nRd02, nRd12,
     nRd22, nRd32);
NR4XB1 I206 ( net053, cds_globals.vdd_, cds_globals.gnd_, net063,
     net016, net057, net054);
NR4XB1 I202 ( net055, cds_globals.vdd_, cds_globals.gnd_, nRd121,
     nRd131, nRd141, nRd151);
NR4XB1 I200 ( net058, cds_globals.vdd_, cds_globals.gnd_, nRd81, nRd91,
     nRd101, nRd111);
NR4XB1 I194 ( net061, cds_globals.vdd_, cds_globals.gnd_, nRd41, nRd51,
     nRd61, nRd71);
NR4XB1 I192 ( net064, cds_globals.vdd_, cds_globals.gnd_, nRd01, nRd11,
     nRd21, nRd31);
NR4XB1 I188 ( net066, cds_globals.vdd_, cds_globals.gnd_, net026,
     net018, net070, net067);
NR4XB1 I184 ( net068, cds_globals.vdd_, cds_globals.gnd_, nRd120,
     nRd130, nRd140, nRd150);
NR4XB1 I182 ( net071, cds_globals.vdd_, cds_globals.gnd_, nRd80, nRd90,
     nRd100, nRd110);
NR4XB1 I177 ( net074, cds_globals.vdd_, cds_globals.gnd_, nRd40, nRd50,
     nRd60, nRd70);
NR4XB1 I171 ( net078, cds_globals.vdd_, cds_globals.gnd_, nRd00, nRd10,
     nRd20, nRd30);
NR4XB1 I148 ( net01, cds_globals.vdd_, cds_globals.gnd_, Rval0, Rval1,
     Rval2, Rval3);
INVXB1 I241 ( Rval3, cds_globals.vdd_, cds_globals.gnd_, net027);
INVXB1 I240 ( net028, cds_globals.vdd_, cds_globals.gnd_, net029);
INVXB1 I233 ( net011, cds_globals.vdd_, cds_globals.gnd_, net032);
INVXB1 I232 ( net012, cds_globals.vdd_, cds_globals.gnd_, net035);
INVXB1 I225 ( net037, cds_globals.vdd_, cds_globals.gnd_, net038);
INVXB1 I223 ( Rval2, cds_globals.vdd_, cds_globals.gnd_, net040);
INVXB1 I222 ( net041, cds_globals.vdd_, cds_globals.gnd_, net042);
INVXB1 I215 ( net013, cds_globals.vdd_, cds_globals.gnd_, net045);
INVXB1 I214 ( net047, cds_globals.vdd_, cds_globals.gnd_, net048);
INVXB1 I207 ( net022, cds_globals.vdd_, cds_globals.gnd_, net051);
INVXB1 I205 ( Rval1, cds_globals.vdd_, cds_globals.gnd_, net053);
INVXB1 I204 ( net054, cds_globals.vdd_, cds_globals.gnd_, net055);
INVXB1 I197 ( net057, cds_globals.vdd_, cds_globals.gnd_, net058);
INVXB1 I196 ( net016, cds_globals.vdd_, cds_globals.gnd_, net061);
INVXB1 I189 ( net063, cds_globals.vdd_, cds_globals.gnd_, net064);
INVXB1 I187 ( Rval0, cds_globals.vdd_, cds_globals.gnd_, net066);
INVXB1 I186 ( net067, cds_globals.vdd_, cds_globals.gnd_, net068);
INVXB1 I179 ( net070, cds_globals.vdd_, cds_globals.gnd_, net071);
INVXB1 I175 ( net018, cds_globals.vdd_, cds_globals.gnd_, net074);
INVXB1 I172 ( net026, cds_globals.vdd_, cds_globals.gnd_, net078);
INVXB1 I149 ( Rval, cds_globals.vdd_, cds_globals.gnd_, net01);

endmodule


// Library - XB16TSMC65, Cell - ZZFBCP, View - schematic
// LAST TIME SAVED: May  8 15:13:02 2023
// NETLIST TIME: May 12 11:49:58 2023
`timescale 1ns / 1ns

module ZZFBCP ( NR00, NR10, NR20, NR30, NR40, NR50, NR60, NR70, NR80,
     NR90, NR100, NR110, NR120, NR130, NR140, NR150, R00, R10, R20,
     R30, R40, R50, R60, R70, R80, R90, R100, R110, R120, R130, R140,
     R150, VDD, VSS, L00, L10, L20, L30, L40, L50, L60, L70, L80, L90,
     L100, L110, L120, L130, L140, L150, NL00, NL10, NL20, NL30, NL40,
     NL50, NL60, NL70, NL80, NL90, NL100, NL110, NL120, NL130, NL140,
     NL150, NRACK0, NRACK1, NRACK2, NRACK3, NRACK4, NRACK5, NRACK6,
     NRACK7, NRACK8, NRACK9, NRACK10, NRACK11, NRACK12, NRACK13,
     NRACK14, NRACK15, NVAL, NX0, NX1, NX2, NX3, NX4, NX5, NX6, NX7,
     NX8, NX9, NX10, NX11, NX12, NX13, NX14, NX15, NX16, NX17, NX18,
     NX19, NX20, NX21, NX22, NX23, NX24, NX25, NX26, NX27, NX28, NX29,
     NX30, NX31, NX32, NX33, NX34, NX35, NX36, NX37, NX38, NX39, NX40,
     NX41, NX42, NX43, NX44, NX45, NX46, NX47, NX48, NX49, NX50, NX51,
     NX52, NX53, NX54, NX55, NX56, NX57, NX58, NX59, NX60, NX61, NX62,
     NX63, NX64, NX65, NX66, NX67, NX68, NX69, NX70, NX71, NX72, NX73,
     NX74, NX75, NX76, NX77, NX78, NX79, NX80, NX81, NX82, NX83, NX84,
     NX85, NX86, NX87, NX88, NX89, NX90, NX91, NX92, NX93, NX94, NX95,
     NX96, NX97, NX98, NX99, NX100, NX101, NX102, NX103, NX104, NX105,
     NX106, NX107, NX108, NX109, NX110, NX111, NX112, NX113, NX114,
     NX115, NX116, NX117, NX118, NX119, NX120, NX121, NX122, NX123,
     NX124, NX125, NX126, NX127, NX128, NX129, NX130, NX131, NX132,
     NX133, NX134, NX135, NX136, NX137, NX138, NX139, NX140, NX141,
     NX142, NX143, NX144, NX145, NX146, NX147, NX148, NX149, NX150,
     NX151, NX152, NX153, NX154, NX155, NX156, NX157, NX158, NX159,
     NX160, NX161, NX162, NX163, NX164, NX165, NX166, NX167, NX168,
     NX169, NX170, NX171, NX172, NX173, NX174, NX175, NX176, NX177,
     NX178, NX179, NX180, NX181, NX182, NX183, NX184, NX185, NX186,
     NX187, NX188, NX189, NX190, NX191, NX192, NX193, NX194, NX195,
     NX196, NX197, NX198, NX199, NX200, NX201, NX202, NX203, NX204,
     NX205, NX206, NX207, NX208, NX209, NX210, NX211, NX212, NX213,
     NX214, NX215, NX216, NX217, NX218, NX219, NX220, NX221, NX222,
     NX223, NX224, NX225, NX226, NX227, NX228, NX229, NX230, NX231,
     NX232, NX233, NX234, NX235, NX236, NX237, NX238, NX239, NX240,
     NX241, NX242, NX243, NX244, NX245, NX246, NX247, NX248, NX249,
     NX250, NX251, NX252, NX253, NX254, NX255, RACK0, RACK1, RACK2,
     RACK3, RACK4, RACK5, RACK6, RACK7, RACK8, RACK9, RACK10, RACK11,
     RACK12, RACK13, RACK14, RACK15, X0, X1, X2, X3, X4, X5, X6, X7,
     X8, X9, X10, X11, X12, X13, X14, X15, X16, X17, X18, X19, X20,
     X21, X22, X23, X24, X25, X26, X27, X28, X29, X30, X31, X32, X33,
     X34, X35, X36, X37, X38, X39, X40, X41, X42, X43, X44, X45, X46,
     X47, X48, X49, X50, X51, X52, X53, X54, X55, X56, X57, X58, X59,
     X60, X61, X62, X63, X64, X65, X66, X67, X68, X69, X70, X71, X72,
     X73, X74, X75, X76, X77, X78, X79, X80, X81, X82, X83, X84, X85,
     X86, X87, X88, X89, X90, X91, X92, X93, X94, X95, X96, X97, X98,
     X99, X100, X101, X102, X103, X104, X105, X106, X107, X108, X109,
     X110, X111, X112, X113, X114, X115, X116, X117, X118, X119, X120,
     X121, X122, X123, X124, X125, X126, X127, X128, X129, X130, X131,
     X132, X133, X134, X135, X136, X137, X138, X139, X140, X141, X142,
     X143, X144, X145, X146, X147, X148, X149, X150, X151, X152, X153,
     X154, X155, X156, X157, X158, X159, X160, X161, X162, X163, X164,
     X165, X166, X167, X168, X169, X170, X171, X172, X173, X174, X175,
     X176, X177, X178, X179, X180, X181, X182, X183, X184, X185, X186,
     X187, X188, X189, X190, X191, X192, X193, X194, X195, X196, X197,
     X198, X199, X200, X201, X202, X203, X204, X205, X206, X207, X208,
     X209, X210, X211, X212, X213, X214, X215, X216, X217, X218, X219,
     X220, X221, X222, X223, X224, X225, X226, X227, X228, X229, X230,
     X231, X232, X233, X234, X235, X236, X237, X238, X239, X240, X241,
     X242, X243, X244, X245, X246, X247, X248, X249, X250, X251, X252,
     X253, X254, X255 );

inout  NR00, NR10, NR20, NR30, NR40, NR50, NR60, NR70, NR80, NR90,
     NR100, NR110, NR120, NR130, NR140, NR150, R00, R10, R20, R30, R40,
     R50, R60, R70, R80, R90, R100, R110, R120, R130, R140, R150, VDD,
     VSS;

input  L00, L10, L20, L30, L40, L50, L60, L70, L80, L90, L100, L110,
     L120, L130, L140, L150, NL00, NL10, NL20, NL30, NL40, NL50, NL60,
     NL70, NL80, NL90, NL100, NL110, NL120, NL130, NL140, NL150,
     NRACK0, NRACK1, NRACK2, NRACK3, NRACK4, NRACK5, NRACK6, NRACK7,
     NRACK8, NRACK9, NRACK10, NRACK11, NRACK12, NRACK13, NRACK14,
     NRACK15, NVAL, NX0, NX1, NX2, NX3, NX4, NX5, NX6, NX7, NX8, NX9,
     NX10, NX11, NX12, NX13, NX14, NX15, NX16, NX17, NX18, NX19, NX20,
     NX21, NX22, NX23, NX24, NX25, NX26, NX27, NX28, NX29, NX30, NX31,
     NX32, NX33, NX34, NX35, NX36, NX37, NX38, NX39, NX40, NX41, NX42,
     NX43, NX44, NX45, NX46, NX47, NX48, NX49, NX50, NX51, NX52, NX53,
     NX54, NX55, NX56, NX57, NX58, NX59, NX60, NX61, NX62, NX63, NX64,
     NX65, NX66, NX67, NX68, NX69, NX70, NX71, NX72, NX73, NX74, NX75,
     NX76, NX77, NX78, NX79, NX80, NX81, NX82, NX83, NX84, NX85, NX86,
     NX87, NX88, NX89, NX90, NX91, NX92, NX93, NX94, NX95, NX96, NX97,
     NX98, NX99, NX100, NX101, NX102, NX103, NX104, NX105, NX106,
     NX107, NX108, NX109, NX110, NX111, NX112, NX113, NX114, NX115,
     NX116, NX117, NX118, NX119, NX120, NX121, NX122, NX123, NX124,
     NX125, NX126, NX127, NX128, NX129, NX130, NX131, NX132, NX133,
     NX134, NX135, NX136, NX137, NX138, NX139, NX140, NX141, NX142,
     NX143, NX144, NX145, NX146, NX147, NX148, NX149, NX150, NX151,
     NX152, NX153, NX154, NX155, NX156, NX157, NX158, NX159, NX160,
     NX161, NX162, NX163, NX164, NX165, NX166, NX167, NX168, NX169,
     NX170, NX171, NX172, NX173, NX174, NX175, NX176, NX177, NX178,
     NX179, NX180, NX181, NX182, NX183, NX184, NX185, NX186, NX187,
     NX188, NX189, NX190, NX191, NX192, NX193, NX194, NX195, NX196,
     NX197, NX198, NX199, NX200, NX201, NX202, NX203, NX204, NX205,
     NX206, NX207, NX208, NX209, NX210, NX211, NX212, NX213, NX214,
     NX215, NX216, NX217, NX218, NX219, NX220, NX221, NX222, NX223,
     NX224, NX225, NX226, NX227, NX228, NX229, NX230, NX231, NX232,
     NX233, NX234, NX235, NX236, NX237, NX238, NX239, NX240, NX241,
     NX242, NX243, NX244, NX245, NX246, NX247, NX248, NX249, NX250,
     NX251, NX252, NX253, NX254, NX255, RACK0, RACK1, RACK2, RACK3,
     RACK4, RACK5, RACK6, RACK7, RACK8, RACK9, RACK10, RACK11, RACK12,
     RACK13, RACK14, RACK15, X0, X1, X2, X3, X4, X5, X6, X7, X8, X9,
     X10, X11, X12, X13, X14, X15, X16, X17, X18, X19, X20, X21, X22,
     X23, X24, X25, X26, X27, X28, X29, X30, X31, X32, X33, X34, X35,
     X36, X37, X38, X39, X40, X41, X42, X43, X44, X45, X46, X47, X48,
     X49, X50, X51, X52, X53, X54, X55, X56, X57, X58, X59, X60, X61,
     X62, X63, X64, X65, X66, X67, X68, X69, X70, X71, X72, X73, X74,
     X75, X76, X77, X78, X79, X80, X81, X82, X83, X84, X85, X86, X87,
     X88, X89, X90, X91, X92, X93, X94, X95, X96, X97, X98, X99, X100,
     X101, X102, X103, X104, X105, X106, X107, X108, X109, X110, X111,
     X112, X113, X114, X115, X116, X117, X118, X119, X120, X121, X122,
     X123, X124, X125, X126, X127, X128, X129, X130, X131, X132, X133,
     X134, X135, X136, X137, X138, X139, X140, X141, X142, X143, X144,
     X145, X146, X147, X148, X149, X150, X151, X152, X153, X154, X155,
     X156, X157, X158, X159, X160, X161, X162, X163, X164, X165, X166,
     X167, X168, X169, X170, X171, X172, X173, X174, X175, X176, X177,
     X178, X179, X180, X181, X182, X183, X184, X185, X186, X187, X188,
     X189, X190, X191, X192, X193, X194, X195, X196, X197, X198, X199,
     X200, X201, X202, X203, X204, X205, X206, X207, X208, X209, X210,
     X211, X212, X213, X214, X215, X216, X217, X218, X219, X220, X221,
     X222, X223, X224, X225, X226, X227, X228, X229, X230, X231, X232,
     X233, X234, X235, X236, X237, X238, X239, X240, X241, X242, X243,
     X244, X245, X246, X247, X248, X249, X250, X251, X252, X253, X254,
     X255;


specify
    specparam CDS_LIBNAME  = "XB16TSMC65";
    specparam CDS_CELLNAME = "ZZFBCP";
    specparam CDS_VIEWNAME = "schematic";
endspecify

CLSAXB1 I285 ( NR40, R40, VDD, VSS, L100, NL100, NRACK4, NVAL, NX164,
     RACK4, X164);
CLSAXB1 I284 ( NR20, R20, VDD, VSS, L100, NL100, NRACK2, NVAL, NX162,
     RACK2, X162);
CLSAXB1 I283 ( NR30, R30, VDD, VSS, L100, NL100, NRACK3, NVAL, NX163,
     RACK3, X163);
CLSAXB1 I282 ( NR00, R00, VDD, VSS, L100, NL100, NRACK0, NVAL, NX160,
     RACK0, X160);
CLSAXB1 I281 ( NR10, R10, VDD, VSS, L100, NL100, NRACK1, NVAL, NX161,
     RACK1, X161);
CLSAXB1 I280 ( NR10, R10, VDD, VSS, L110, NL110, NRACK1, NVAL, NX177,
     RACK1, X177);
CLSAXB1 I279 ( NR20, R20, VDD, VSS, L110, NL110, NRACK2, NVAL, NX178,
     RACK2, X178);
CLSAXB1 I278 ( NR30, R30, VDD, VSS, L110, NL110, NRACK3, NVAL, NX179,
     RACK3, X179);
CLSAXB1 I277 ( NR40, R40, VDD, VSS, L110, NL110, NRACK4, NVAL, NX180,
     RACK4, X180);
CLSAXB1 I276 ( NR40, R40, VDD, VSS, L120, NL120, NRACK4, NVAL, NX196,
     RACK4, X196);
CLSAXB1 I275 ( NR30, R30, VDD, VSS, L120, NL120, NRACK3, NVAL, NX195,
     RACK3, X195);
CLSAXB1 I274 ( NR20, R20, VDD, VSS, L120, NL120, NRACK2, NVAL, NX194,
     RACK2, X194);
CLSAXB1 I273 ( NR10, R10, VDD, VSS, L120, NL120, NRACK1, NVAL, NX193,
     RACK1, X193);
CLSAXB1 I272 ( NR00, R00, VDD, VSS, L120, NL120, NRACK0, NVAL, NX192,
     RACK0, X192);
CLSAXB1 I271 ( NR00, R00, VDD, VSS, L130, NL130, NRACK0, NVAL, NX208,
     RACK0, X208);
CLSAXB1 I270 ( NR10, R10, VDD, VSS, L130, NL130, NRACK1, NVAL, NX209,
     RACK1, X209);
CLSAXB1 I269 ( NR20, R20, VDD, VSS, L130, NL130, NRACK2, NVAL, NX210,
     RACK2, X210);
CLSAXB1 I268 ( NR30, R30, VDD, VSS, L130, NL130, NRACK3, NVAL, NX211,
     RACK3, X211);
CLSAXB1 I267 ( NR40, R40, VDD, VSS, L130, NL130, NRACK4, NVAL, NX212,
     RACK4, X212);
CLSAXB1 I266 ( NR40, R40, VDD, VSS, L140, NL140, NRACK4, NVAL, NX228,
     RACK4, X228);
CLSAXB1 I265 ( NR30, R30, VDD, VSS, L140, NL140, NRACK3, NVAL, NX227,
     RACK3, X227);
CLSAXB1 I264 ( NR20, R20, VDD, VSS, L140, NL140, NRACK2, NVAL, NX226,
     RACK2, X226);
CLSAXB1 I263 ( NR00, R00, VDD, VSS, L140, NL140, NRACK0, NVAL, NX224,
     RACK0, X224);
CLSAXB1 I262 ( NR10, R10, VDD, VSS, L140, NL140, NRACK1, NVAL, NX225,
     RACK1, X225);
CLSAXB1 I261 ( NR40, R40, VDD, VSS, L150, NL150, NRACK4, NVAL, NX244,
     RACK4, X244);
CLSAXB1 I260 ( NR20, R20, VDD, VSS, L150, NL150, NRACK2, NVAL, NX242,
     RACK2, X242);
CLSAXB1 I259 ( NR30, R30, VDD, VSS, L150, NL150, NRACK3, NVAL, NX243,
     RACK3, X243);
CLSAXB1 I258 ( NR00, R00, VDD, VSS, L150, NL150, NRACK0, NVAL, NX240,
     RACK0, X240);
CLSAXB1 I257 ( NR10, R10, VDD, VSS, L150, NL150, NRACK1, NVAL, NX241,
     RACK1, X241);
CLSAXB1 I256 ( NR00, R00, VDD, VSS, L110, NL110, NRACK0, NVAL, NX176,
     RACK0, X176);
CLSAXB1 I255 ( NR150, R150, VDD, VSS, L110, NL110, NRACK15, NVAL,
     NX191, RACK15, X191);
CLSAXB1 I254 ( NR150, R150, VDD, VSS, L120, NL120, NRACK15, NVAL,
     NX207, RACK15, X207);
CLSAXB1 I253 ( NR150, R150, VDD, VSS, L130, NL130, NRACK15, NVAL,
     NX223, RACK15, X223);
CLSAXB1 I252 ( NR150, R150, VDD, VSS, L140, NL140, NRACK15, NVAL,
     NX239, RACK15, X239);
CLSAXB1 I251 ( NR150, R150, VDD, VSS, L150, NL150, NRACK15, NVAL,
     NX255, RACK15, X255);
CLSAXB1 I250 ( NR110, R110, VDD, VSS, L110, NL110, NRACK11, NVAL,
     NX187, RACK11, X187);
CLSAXB1 I249 ( NR120, R120, VDD, VSS, L110, NL110, NRACK12, NVAL,
     NX188, RACK12, X188);
CLSAXB1 I248 ( NR130, R130, VDD, VSS, L110, NL110, NRACK13, NVAL,
     NX189, RACK13, X189);
CLSAXB1 I247 ( NR140, R140, VDD, VSS, L110, NL110, NRACK14, NVAL,
     NX190, RACK14, X190);
CLSAXB1 I246 ( NR140, R140, VDD, VSS, L120, NL120, NRACK14, NVAL,
     NX206, RACK14, X206);
CLSAXB1 I245 ( NR130, R130, VDD, VSS, L120, NL120, NRACK13, NVAL,
     NX205, RACK13, X205);
CLSAXB1 I244 ( NR120, R120, VDD, VSS, L120, NL120, NRACK12, NVAL,
     NX204, RACK12, X204);
CLSAXB1 I243 ( NR110, R110, VDD, VSS, L120, NL120, NRACK11, NVAL,
     NX203, RACK11, X203);
CLSAXB1 I242 ( NR100, R100, VDD, VSS, L120, NL120, NRACK10, NVAL,
     NX202, RACK10, X202);
CLSAXB1 I241 ( NR100, R100, VDD, VSS, L130, NL130, NRACK10, NVAL,
     NX218, RACK10, X218);
CLSAXB1 I240 ( NR110, R110, VDD, VSS, L130, NL130, NRACK11, NVAL,
     NX219, RACK11, X219);
CLSAXB1 I239 ( NR120, R120, VDD, VSS, L130, NL130, NRACK12, NVAL,
     NX220, RACK12, X220);
CLSAXB1 I238 ( NR130, R130, VDD, VSS, L130, NL130, NRACK13, NVAL,
     NX221, RACK13, X221);
CLSAXB1 I237 ( NR140, R140, VDD, VSS, L130, NL130, NRACK14, NVAL,
     NX222, RACK14, X222);
CLSAXB1 I236 ( NR140, R140, VDD, VSS, L140, NL140, NRACK14, NVAL,
     NX238, RACK14, X238);
CLSAXB1 I235 ( NR130, R130, VDD, VSS, L140, NL140, NRACK13, NVAL,
     NX237, RACK13, X237);
CLSAXB1 I234 ( NR120, R120, VDD, VSS, L140, NL140, NRACK12, NVAL,
     NX236, RACK12, X236);
CLSAXB1 I233 ( NR100, R100, VDD, VSS, L140, NL140, NRACK10, NVAL,
     NX234, RACK10, X234);
CLSAXB1 I232 ( NR110, R110, VDD, VSS, L140, NL140, NRACK11, NVAL,
     NX235, RACK11, X235);
CLSAXB1 I231 ( NR140, R140, VDD, VSS, L150, NL150, NRACK14, NVAL,
     NX254, RACK14, X254);
CLSAXB1 I230 ( NR120, R120, VDD, VSS, L150, NL150, NRACK12, NVAL,
     NX252, RACK12, X252);
CLSAXB1 I229 ( NR130, R130, VDD, VSS, L150, NL150, NRACK13, NVAL,
     NX253, RACK13, X253);
CLSAXB1 I228 ( NR100, R100, VDD, VSS, L150, NL150, NRACK10, NVAL,
     NX250, RACK10, X250);
CLSAXB1 I227 ( NR110, R110, VDD, VSS, L150, NL150, NRACK11, NVAL,
     NX251, RACK11, X251);
CLSAXB1 I226 ( NR100, R100, VDD, VSS, L110, NL110, NRACK10, NVAL,
     NX186, RACK10, X186);
CLSAXB1 I225 ( NR60, R60, VDD, VSS, L110, NL110, NRACK6, NVAL, NX182,
     RACK6, X182);
CLSAXB1 I224 ( NR70, R70, VDD, VSS, L110, NL110, NRACK7, NVAL, NX183,
     RACK7, X183);
CLSAXB1 I223 ( NR80, R80, VDD, VSS, L110, NL110, NRACK8, NVAL, NX184,
     RACK8, X184);
CLSAXB1 I222 ( NR90, R90, VDD, VSS, L110, NL110, NRACK9, NVAL, NX185,
     RACK9, X185);
CLSAXB1 I221 ( NR90, R90, VDD, VSS, L120, NL120, NRACK9, NVAL, NX201,
     RACK9, X201);
CLSAXB1 I220 ( NR80, R80, VDD, VSS, L120, NL120, NRACK8, NVAL, NX200,
     RACK8, X200);
CLSAXB1 I219 ( NR70, R70, VDD, VSS, L120, NL120, NRACK7, NVAL, NX199,
     RACK7, X199);
CLSAXB1 I218 ( NR60, R60, VDD, VSS, L120, NL120, NRACK6, NVAL, NX198,
     RACK6, X198);
CLSAXB1 I217 ( NR50, R50, VDD, VSS, L120, NL120, NRACK5, NVAL, NX197,
     RACK5, X197);
CLSAXB1 I216 ( NR50, R50, VDD, VSS, L130, NL130, NRACK5, NVAL, NX213,
     RACK5, X213);
CLSAXB1 I215 ( NR60, R60, VDD, VSS, L130, NL130, NRACK6, NVAL, NX214,
     RACK6, X214);
CLSAXB1 I214 ( NR70, R70, VDD, VSS, L130, NL130, NRACK7, NVAL, NX215,
     RACK7, X215);
CLSAXB1 I213 ( NR80, R80, VDD, VSS, L130, NL130, NRACK8, NVAL, NX216,
     RACK8, X216);
CLSAXB1 I212 ( NR90, R90, VDD, VSS, L130, NL130, NRACK9, NVAL, NX217,
     RACK9, X217);
CLSAXB1 I211 ( NR90, R90, VDD, VSS, L140, NL140, NRACK9, NVAL, NX233,
     RACK9, X233);
CLSAXB1 I210 ( NR80, R80, VDD, VSS, L140, NL140, NRACK8, NVAL, NX232,
     RACK8, X232);
CLSAXB1 I209 ( NR70, R70, VDD, VSS, L140, NL140, NRACK7, NVAL, NX231,
     RACK7, X231);
CLSAXB1 I208 ( NR50, R50, VDD, VSS, L140, NL140, NRACK5, NVAL, NX229,
     RACK5, X229);
CLSAXB1 I207 ( NR60, R60, VDD, VSS, L140, NL140, NRACK6, NVAL, NX230,
     RACK6, X230);
CLSAXB1 I206 ( NR90, R90, VDD, VSS, L150, NL150, NRACK9, NVAL, NX249,
     RACK9, X249);
CLSAXB1 I205 ( NR70, R70, VDD, VSS, L150, NL150, NRACK7, NVAL, NX247,
     RACK7, X247);
CLSAXB1 I204 ( NR80, R80, VDD, VSS, L150, NL150, NRACK8, NVAL, NX248,
     RACK8, X248);
CLSAXB1 I203 ( NR50, R50, VDD, VSS, L150, NL150, NRACK5, NVAL, NX245,
     RACK5, X245);
CLSAXB1 I202 ( NR60, R60, VDD, VSS, L150, NL150, NRACK6, NVAL, NX246,
     RACK6, X246);
CLSAXB1 I201 ( NR50, R50, VDD, VSS, L110, NL110, NRACK5, NVAL, NX181,
     RACK5, X181);
CLSAXB1 I200 ( NR150, R150, VDD, VSS, L100, NL100, NRACK15, NVAL,
     NX175, RACK15, X175);
CLSAXB1 I199 ( NR140, R140, VDD, VSS, L100, NL100, NRACK14, NVAL,
     NX174, RACK14, X174);
CLSAXB1 I198 ( NR120, R120, VDD, VSS, L100, NL100, NRACK12, NVAL,
     NX172, RACK12, X172);
CLSAXB1 I197 ( NR130, R130, VDD, VSS, L100, NL100, NRACK13, NVAL,
     NX173, RACK13, X173);
CLSAXB1 I196 ( NR100, R100, VDD, VSS, L100, NL100, NRACK10, NVAL,
     NX170, RACK10, X170);
CLSAXB1 I195 ( NR110, R110, VDD, VSS, L100, NL100, NRACK11, NVAL,
     NX171, RACK11, X171);
CLSAXB1 I194 ( NR90, R90, VDD, VSS, L100, NL100, NRACK9, NVAL, NX169,
     RACK9, X169);
CLSAXB1 I193 ( NR70, R70, VDD, VSS, L100, NL100, NRACK7, NVAL, NX167,
     RACK7, X167);
CLSAXB1 I192 ( NR80, R80, VDD, VSS, L100, NL100, NRACK8, NVAL, NX168,
     RACK8, X168);
CLSAXB1 I191 ( NR50, R50, VDD, VSS, L100, NL100, NRACK5, NVAL, NX165,
     RACK5, X165);
CLSAXB1 I190 ( NR60, R60, VDD, VSS, L100, NL100, NRACK6, NVAL, NX166,
     RACK6, X166);
CLSAXB1 I189 ( NR10, R10, VDD, VSS, L50, NL50, NRACK1, NVAL, NX81,
     RACK1, X81);
CLSAXB1 I188 ( NR20, R20, VDD, VSS, L50, NL50, NRACK2, NVAL, NX82,
     RACK2, X82);
CLSAXB1 I187 ( NR30, R30, VDD, VSS, L50, NL50, NRACK3, NVAL, NX83,
     RACK3, X83);
CLSAXB1 I186 ( NR40, R40, VDD, VSS, L50, NL50, NRACK4, NVAL, NX84,
     RACK4, X84);
CLSAXB1 I185 ( NR40, R40, VDD, VSS, L60, NL60, NRACK4, NVAL, NX100,
     RACK4, X100);
CLSAXB1 I184 ( NR30, R30, VDD, VSS, L60, NL60, NRACK3, NVAL, NX99,
     RACK3, X99);
CLSAXB1 I183 ( NR20, R20, VDD, VSS, L60, NL60, NRACK2, NVAL, NX98,
     RACK2, X98);
CLSAXB1 I182 ( NR10, R10, VDD, VSS, L60, NL60, NRACK1, NVAL, NX97,
     RACK1, X97);
CLSAXB1 I181 ( NR00, R00, VDD, VSS, L60, NL60, NRACK0, NVAL, NX96,
     RACK0, X96);
CLSAXB1 I180 ( NR00, R00, VDD, VSS, L70, NL70, NRACK0, NVAL, NX112,
     RACK0, X112);
CLSAXB1 I179 ( NR10, R10, VDD, VSS, L70, NL70, NRACK1, NVAL, NX113,
     RACK1, X113);
CLSAXB1 I178 ( NR20, R20, VDD, VSS, L70, NL70, NRACK2, NVAL, NX114,
     RACK2, X114);
CLSAXB1 I177 ( NR30, R30, VDD, VSS, L70, NL70, NRACK3, NVAL, NX115,
     RACK3, X115);
CLSAXB1 I176 ( NR40, R40, VDD, VSS, L70, NL70, NRACK4, NVAL, NX116,
     RACK4, X116);
CLSAXB1 I175 ( NR40, R40, VDD, VSS, L80, NL80, NRACK4, NVAL, NX132,
     RACK4, X132);
CLSAXB1 I174 ( NR30, R30, VDD, VSS, L80, NL80, NRACK3, NVAL, NX131,
     RACK3, X131);
CLSAXB1 I173 ( NR20, R20, VDD, VSS, L80, NL80, NRACK2, NVAL, NX130,
     RACK2, X130);
CLSAXB1 I172 ( NR00, R00, VDD, VSS, L80, NL80, NRACK0, NVAL, NX128,
     RACK0, X128);
CLSAXB1 I171 ( NR10, R10, VDD, VSS, L80, NL80, NRACK1, NVAL, NX129,
     RACK1, X129);
CLSAXB1 I170 ( NR40, R40, VDD, VSS, L90, NL90, NRACK4, NVAL, NX148,
     RACK4, X148);
CLSAXB1 I169 ( NR20, R20, VDD, VSS, L90, NL90, NRACK2, NVAL, NX146,
     RACK2, X146);
CLSAXB1 I168 ( NR30, R30, VDD, VSS, L90, NL90, NRACK3, NVAL, NX147,
     RACK3, X147);
CLSAXB1 I167 ( NR00, R00, VDD, VSS, L90, NL90, NRACK0, NVAL, NX144,
     RACK0, X144);
CLSAXB1 I166 ( NR10, R10, VDD, VSS, L90, NL90, NRACK1, NVAL, NX145,
     RACK1, X145);
CLSAXB1 I165 ( NR00, R00, VDD, VSS, L50, NL50, NRACK0, NVAL, NX80,
     RACK0, X80);
CLSAXB1 I164 ( NR150, R150, VDD, VSS, L50, NL50, NRACK15, NVAL, NX95,
     RACK15, X95);
CLSAXB1 I163 ( NR150, R150, VDD, VSS, L60, NL60, NRACK15, NVAL, NX111,
     RACK15, X111);
CLSAXB1 I162 ( NR150, R150, VDD, VSS, L70, NL70, NRACK15, NVAL, NX127,
     RACK15, X127);
CLSAXB1 I161 ( NR150, R150, VDD, VSS, L80, NL80, NRACK15, NVAL, NX143,
     RACK15, X143);
CLSAXB1 I160 ( NR150, R150, VDD, VSS, L90, NL90, NRACK15, NVAL, NX159,
     RACK15, X159);
CLSAXB1 I159 ( NR110, R110, VDD, VSS, L50, NL50, NRACK11, NVAL, NX91,
     RACK11, X91);
CLSAXB1 I158 ( NR120, R120, VDD, VSS, L50, NL50, NRACK12, NVAL, NX92,
     RACK12, X92);
CLSAXB1 I157 ( NR130, R130, VDD, VSS, L50, NL50, NRACK13, NVAL, NX93,
     RACK13, X93);
CLSAXB1 I156 ( NR140, R140, VDD, VSS, L50, NL50, NRACK14, NVAL, NX94,
     RACK14, X94);
CLSAXB1 I155 ( NR140, R140, VDD, VSS, L60, NL60, NRACK14, NVAL, NX110,
     RACK14, X110);
CLSAXB1 I154 ( NR130, R130, VDD, VSS, L60, NL60, NRACK13, NVAL, NX109,
     RACK13, X109);
CLSAXB1 I153 ( NR120, R120, VDD, VSS, L60, NL60, NRACK12, NVAL, NX108,
     RACK12, X108);
CLSAXB1 I152 ( NR110, R110, VDD, VSS, L60, NL60, NRACK11, NVAL, NX107,
     RACK11, X107);
CLSAXB1 I151 ( NR100, R100, VDD, VSS, L60, NL60, NRACK10, NVAL, NX106,
     RACK10, X106);
CLSAXB1 I150 ( NR100, R100, VDD, VSS, L70, NL70, NRACK10, NVAL, NX122,
     RACK10, X122);
CLSAXB1 I149 ( NR110, R110, VDD, VSS, L70, NL70, NRACK11, NVAL, NX123,
     RACK11, X123);
CLSAXB1 I148 ( NR120, R120, VDD, VSS, L70, NL70, NRACK12, NVAL, NX124,
     RACK12, X124);
CLSAXB1 I147 ( NR130, R130, VDD, VSS, L70, NL70, NRACK13, NVAL, NX125,
     RACK13, X125);
CLSAXB1 I146 ( NR140, R140, VDD, VSS, L70, NL70, NRACK14, NVAL, NX126,
     RACK14, X126);
CLSAXB1 I145 ( NR140, R140, VDD, VSS, L80, NL80, NRACK14, NVAL, NX142,
     RACK14, X142);
CLSAXB1 I144 ( NR130, R130, VDD, VSS, L80, NL80, NRACK13, NVAL, NX141,
     RACK13, X141);
CLSAXB1 I143 ( NR120, R120, VDD, VSS, L80, NL80, NRACK12, NVAL, NX140,
     RACK12, X140);
CLSAXB1 I142 ( NR100, R100, VDD, VSS, L80, NL80, NRACK10, NVAL, NX138,
     RACK10, X138);
CLSAXB1 I141 ( NR110, R110, VDD, VSS, L80, NL80, NRACK11, NVAL, NX139,
     RACK11, X139);
CLSAXB1 I140 ( NR140, R140, VDD, VSS, L90, NL90, NRACK14, NVAL, NX158,
     RACK14, X158);
CLSAXB1 I139 ( NR120, R120, VDD, VSS, L90, NL90, NRACK12, NVAL, NX156,
     RACK12, X156);
CLSAXB1 I138 ( NR130, R130, VDD, VSS, L90, NL90, NRACK13, NVAL, NX157,
     RACK13, X157);
CLSAXB1 I137 ( NR100, R100, VDD, VSS, L90, NL90, NRACK10, NVAL, NX154,
     RACK10, X154);
CLSAXB1 I136 ( NR110, R110, VDD, VSS, L90, NL90, NRACK11, NVAL, NX155,
     RACK11, X155);
CLSAXB1 I135 ( NR100, R100, VDD, VSS, L50, NL50, NRACK10, NVAL, NX90,
     RACK10, X90);
CLSAXB1 I134 ( NR60, R60, VDD, VSS, L50, NL50, NRACK6, NVAL, NX86,
     RACK6, X86);
CLSAXB1 I133 ( NR70, R70, VDD, VSS, L50, NL50, NRACK7, NVAL, NX87,
     RACK7, X87);
CLSAXB1 I132 ( NR80, R80, VDD, VSS, L50, NL50, NRACK8, NVAL, NX88,
     RACK8, X88);
CLSAXB1 I131 ( NR90, R90, VDD, VSS, L50, NL50, NRACK9, NVAL, NX89,
     RACK9, X89);
CLSAXB1 I130 ( NR90, R90, VDD, VSS, L60, NL60, NRACK9, NVAL, NX105,
     RACK9, X105);
CLSAXB1 I129 ( NR80, R80, VDD, VSS, L60, NL60, NRACK8, NVAL, NX104,
     RACK8, X104);
CLSAXB1 I128 ( NR70, R70, VDD, VSS, L60, NL60, NRACK7, NVAL, NX103,
     RACK7, X103);
CLSAXB1 I127 ( NR60, R60, VDD, VSS, L60, NL60, NRACK6, NVAL, NX102,
     RACK6, X102);
CLSAXB1 I126 ( NR50, R50, VDD, VSS, L60, NL60, NRACK5, NVAL, NX101,
     RACK5, X101);
CLSAXB1 I125 ( NR50, R50, VDD, VSS, L70, NL70, NRACK5, NVAL, NX117,
     RACK5, X117);
CLSAXB1 I124 ( NR60, R60, VDD, VSS, L70, NL70, NRACK6, NVAL, NX118,
     RACK6, X118);
CLSAXB1 I123 ( NR70, R70, VDD, VSS, L70, NL70, NRACK7, NVAL, NX119,
     RACK7, X119);
CLSAXB1 I122 ( NR80, R80, VDD, VSS, L70, NL70, NRACK8, NVAL, NX120,
     RACK8, X120);
CLSAXB1 I121 ( NR90, R90, VDD, VSS, L70, NL70, NRACK9, NVAL, NX121,
     RACK9, X121);
CLSAXB1 I120 ( NR90, R90, VDD, VSS, L80, NL80, NRACK9, NVAL, NX137,
     RACK9, X137);
CLSAXB1 I119 ( NR80, R80, VDD, VSS, L80, NL80, NRACK8, NVAL, NX136,
     RACK8, X136);
CLSAXB1 I118 ( NR70, R70, VDD, VSS, L80, NL80, NRACK7, NVAL, NX135,
     RACK7, X135);
CLSAXB1 I117 ( NR50, R50, VDD, VSS, L80, NL80, NRACK5, NVAL, NX133,
     RACK5, X133);
CLSAXB1 I116 ( NR60, R60, VDD, VSS, L80, NL80, NRACK6, NVAL, NX134,
     RACK6, X134);
CLSAXB1 I115 ( NR90, R90, VDD, VSS, L90, NL90, NRACK9, NVAL, NX153,
     RACK9, X153);
CLSAXB1 I114 ( NR70, R70, VDD, VSS, L90, NL90, NRACK7, NVAL, NX151,
     RACK7, X151);
CLSAXB1 I113 ( NR80, R80, VDD, VSS, L90, NL90, NRACK8, NVAL, NX152,
     RACK8, X152);
CLSAXB1 I112 ( NR50, R50, VDD, VSS, L90, NL90, NRACK5, NVAL, NX149,
     RACK5, X149);
CLSAXB1 I111 ( NR60, R60, VDD, VSS, L90, NL90, NRACK6, NVAL, NX150,
     RACK6, X150);
CLSAXB1 I110 ( NR50, R50, VDD, VSS, L50, NL50, NRACK5, NVAL, NX85,
     RACK5, X85);
CLSAXB1 I109 ( NR150, R150, VDD, VSS, L00, NL00, NRACK15, NVAL, NX15,
     RACK15, X15);
CLSAXB1 I108 ( NR150, R150, VDD, VSS, L10, NL10, NRACK15, NVAL, NX31,
     RACK15, X31);
CLSAXB1 I107 ( NR150, R150, VDD, VSS, L20, NL20, NRACK15, NVAL, NX47,
     RACK15, X47);
CLSAXB1 I106 ( NR150, R150, VDD, VSS, L30, NL30, NRACK15, NVAL, NX63,
     RACK15, X63);
CLSAXB1 I105 ( NR150, R150, VDD, VSS, L40, NL40, NRACK15, NVAL, NX79,
     RACK15, X79);
CLSAXB1 I104 ( NR110, R110, VDD, VSS, L00, NL00, NRACK11, NVAL, NX11,
     RACK11, X11);
CLSAXB1 I103 ( NR120, R120, VDD, VSS, L00, NL00, NRACK12, NVAL, NX12,
     RACK12, X12);
CLSAXB1 I102 ( NR130, R130, VDD, VSS, L00, NL00, NRACK13, NVAL, NX13,
     RACK13, X13);
CLSAXB1 I101 ( NR140, R140, VDD, VSS, L00, NL00, NRACK14, NVAL, NX14,
     RACK14, X14);
CLSAXB1 I100 ( NR140, R140, VDD, VSS, L10, NL10, NRACK14, NVAL, NX30,
     RACK14, X30);
CLSAXB1 I99 ( NR130, R130, VDD, VSS, L10, NL10, NRACK13, NVAL, NX29,
     RACK13, X29);
CLSAXB1 I98 ( NR120, R120, VDD, VSS, L10, NL10, NRACK12, NVAL, NX28,
     RACK12, X28);
CLSAXB1 I97 ( NR110, R110, VDD, VSS, L10, NL10, NRACK11, NVAL, NX27,
     RACK11, X27);
CLSAXB1 I96 ( NR100, R100, VDD, VSS, L10, NL10, NRACK10, NVAL, NX26,
     RACK10, X26);
CLSAXB1 I95 ( NR100, R100, VDD, VSS, L20, NL20, NRACK10, NVAL, NX42,
     RACK10, X42);
CLSAXB1 I94 ( NR110, R110, VDD, VSS, L20, NL20, NRACK11, NVAL, NX43,
     RACK11, X43);
CLSAXB1 I93 ( NR120, R120, VDD, VSS, L20, NL20, NRACK12, NVAL, NX44,
     RACK12, X44);
CLSAXB1 I92 ( NR130, R130, VDD, VSS, L20, NL20, NRACK13, NVAL, NX45,
     RACK13, X45);
CLSAXB1 I91 ( NR140, R140, VDD, VSS, L20, NL20, NRACK14, NVAL, NX46,
     RACK14, X46);
CLSAXB1 I90 ( NR140, R140, VDD, VSS, L30, NL30, NRACK14, NVAL, NX62,
     RACK14, X62);
CLSAXB1 I89 ( NR130, R130, VDD, VSS, L30, NL30, NRACK13, NVAL, NX61,
     RACK13, X61);
CLSAXB1 I88 ( NR120, R120, VDD, VSS, L30, NL30, NRACK12, NVAL, NX60,
     RACK12, X60);
CLSAXB1 I87 ( NR100, R100, VDD, VSS, L30, NL30, NRACK10, NVAL, NX58,
     RACK10, X58);
CLSAXB1 I86 ( NR110, R110, VDD, VSS, L30, NL30, NRACK11, NVAL, NX59,
     RACK11, X59);
CLSAXB1 I85 ( NR140, R140, VDD, VSS, L40, NL40, NRACK14, NVAL, NX78,
     RACK14, X78);
CLSAXB1 I84 ( NR120, R120, VDD, VSS, L40, NL40, NRACK12, NVAL, NX76,
     RACK12, X76);
CLSAXB1 I83 ( NR130, R130, VDD, VSS, L40, NL40, NRACK13, NVAL, NX77,
     RACK13, X77);
CLSAXB1 I82 ( NR100, R100, VDD, VSS, L40, NL40, NRACK10, NVAL, NX74,
     RACK10, X74);
CLSAXB1 I81 ( NR110, R110, VDD, VSS, L40, NL40, NRACK11, NVAL, NX75,
     RACK11, X75);
CLSAXB1 I80 ( NR100, R100, VDD, VSS, L00, NL00, NRACK10, NVAL, NX10,
     RACK10, X10);
CLSAXB1 I79 ( NR60, R60, VDD, VSS, L00, NL00, NRACK6, NVAL, NX6, RACK6,
     X6);
CLSAXB1 I78 ( NR70, R70, VDD, VSS, L00, NL00, NRACK7, NVAL, NX7, RACK7,
     X7);
CLSAXB1 I77 ( NR80, R80, VDD, VSS, L00, NL00, NRACK8, NVAL, NX8, RACK8,
     X8);
CLSAXB1 I76 ( NR90, R90, VDD, VSS, L00, NL00, NRACK9, NVAL, NX9, RACK9,
     X9);
CLSAXB1 I75 ( NR90, R90, VDD, VSS, L10, NL10, NRACK9, NVAL, NX25,
     RACK9, X25);
CLSAXB1 I74 ( NR80, R80, VDD, VSS, L10, NL10, NRACK8, NVAL, NX24,
     RACK8, X24);
CLSAXB1 I73 ( NR70, R70, VDD, VSS, L10, NL10, NRACK7, NVAL, NX23,
     RACK7, X23);
CLSAXB1 I72 ( NR60, R60, VDD, VSS, L10, NL10, NRACK6, NVAL, NX22,
     RACK6, X22);
CLSAXB1 I71 ( NR50, R50, VDD, VSS, L10, NL10, NRACK5, NVAL, NX21,
     RACK5, X21);
CLSAXB1 I70 ( NR50, R50, VDD, VSS, L20, NL20, NRACK5, NVAL, NX37,
     RACK5, X37);
CLSAXB1 I69 ( NR60, R60, VDD, VSS, L20, NL20, NRACK6, NVAL, NX38,
     RACK6, X38);
CLSAXB1 I68 ( NR70, R70, VDD, VSS, L20, NL20, NRACK7, NVAL, NX39,
     RACK7, X39);
CLSAXB1 I67 ( NR80, R80, VDD, VSS, L20, NL20, NRACK8, NVAL, NX40,
     RACK8, X40);
CLSAXB1 I66 ( NR90, R90, VDD, VSS, L20, NL20, NRACK9, NVAL, NX41,
     RACK9, X41);
CLSAXB1 I65 ( NR90, R90, VDD, VSS, L30, NL30, NRACK9, NVAL, NX57,
     RACK9, X57);
CLSAXB1 I64 ( NR80, R80, VDD, VSS, L30, NL30, NRACK8, NVAL, NX56,
     RACK8, X56);
CLSAXB1 I63 ( NR70, R70, VDD, VSS, L30, NL30, NRACK7, NVAL, NX55,
     RACK7, X55);
CLSAXB1 I62 ( NR50, R50, VDD, VSS, L30, NL30, NRACK5, NVAL, NX53,
     RACK5, X53);
CLSAXB1 I61 ( NR60, R60, VDD, VSS, L30, NL30, NRACK6, NVAL, NX54,
     RACK6, X54);
CLSAXB1 I60 ( NR90, R90, VDD, VSS, L40, NL40, NRACK9, NVAL, NX73,
     RACK9, X73);
CLSAXB1 I59 ( NR70, R70, VDD, VSS, L40, NL40, NRACK7, NVAL, NX71,
     RACK7, X71);
CLSAXB1 I58 ( NR80, R80, VDD, VSS, L40, NL40, NRACK8, NVAL, NX72,
     RACK8, X72);
CLSAXB1 I57 ( NR50, R50, VDD, VSS, L40, NL40, NRACK5, NVAL, NX69,
     RACK5, X69);
CLSAXB1 I56 ( NR60, R60, VDD, VSS, L40, NL40, NRACK6, NVAL, NX70,
     RACK6, X70);
CLSAXB1 I50 ( NR40, R40, VDD, VSS, L40, NL40, NRACK4, NVAL, NX68,
     RACK4, X68);
CLSAXB1 I52 ( NR20, R20, VDD, VSS, L40, NL40, NRACK2, NVAL, NX66,
     RACK2, X66);
CLSAXB1 I51 ( NR30, R30, VDD, VSS, L40, NL40, NRACK3, NVAL, NX67,
     RACK3, X67);
CLSAXB1 I54 ( NR00, R00, VDD, VSS, L40, NL40, NRACK0, NVAL, NX64,
     RACK0, X64);
CLSAXB1 I53 ( NR10, R10, VDD, VSS, L40, NL40, NRACK1, NVAL, NX65,
     RACK1, X65);
CLSAXB1 I45 ( NR40, R40, VDD, VSS, L30, NL30, NRACK4, NVAL, NX52,
     RACK4, X52);
CLSAXB1 I46 ( NR30, R30, VDD, VSS, L30, NL30, NRACK3, NVAL, NX51,
     RACK3, X51);
CLSAXB1 I47 ( NR20, R20, VDD, VSS, L30, NL30, NRACK2, NVAL, NX50,
     RACK2, X50);
CLSAXB1 I31 ( NR10, R10, VDD, VSS, L00, NL00, NRACK1, NVAL, NX1, RACK1,
     X1);
CLSAXB1 I30 ( NR00, R00, VDD, VSS, L00, NL00, NRACK0, NVAL, NX0, RACK0,
     X0);
CLSAXB1 I55 ( NR50, R50, VDD, VSS, L00, NL00, NRACK5, NVAL, NX5, RACK5,
     X5);
CLSAXB1 I39 ( NR40, R40, VDD, VSS, L10, NL10, NRACK4, NVAL, NX20,
     RACK4, X20);
CLSAXB1 I38 ( NR30, R30, VDD, VSS, L10, NL10, NRACK3, NVAL, NX19,
     RACK3, X19);
CLSAXB1 I37 ( NR20, R20, VDD, VSS, L10, NL10, NRACK2, NVAL, NX18,
     RACK2, X18);
CLSAXB1 I36 ( NR10, R10, VDD, VSS, L10, NL10, NRACK1, NVAL, NX17,
     RACK1, X17);
CLSAXB1 I32 ( NR20, R20, VDD, VSS, L00, NL00, NRACK2, NVAL, NX2, RACK2,
     X2);
CLSAXB1 I33 ( NR30, R30, VDD, VSS, L00, NL00, NRACK3, NVAL, NX3, RACK3,
     X3);
CLSAXB1 I34 ( NR40, R40, VDD, VSS, L00, NL00, NRACK4, NVAL, NX4, RACK4,
     X4);
CLSAXB1 I35 ( NR00, R00, VDD, VSS, L10, NL10, NRACK0, NVAL, NX16,
     RACK0, X16);
CLSAXB1 I44 ( NR00, R00, VDD, VSS, L20, NL20, NRACK0, NVAL, NX32,
     RACK0, X32);
CLSAXB1 I43 ( NR10, R10, VDD, VSS, L20, NL20, NRACK1, NVAL, NX33,
     RACK1, X33);
CLSAXB1 I42 ( NR20, R20, VDD, VSS, L20, NL20, NRACK2, NVAL, NX34,
     RACK2, X34);
CLSAXB1 I41 ( NR30, R30, VDD, VSS, L20, NL20, NRACK3, NVAL, NX35,
     RACK3, X35);
CLSAXB1 I40 ( NR40, R40, VDD, VSS, L20, NL20, NRACK4, NVAL, NX36,
     RACK4, X36);
CLSAXB1 I49 ( NR00, R00, VDD, VSS, L30, NL30, NRACK0, NVAL, NX48,
     RACK0, X48);
CLSAXB1 I48 ( NR10, R10, VDD, VSS, L30, NL30, NRACK1, NVAL, NX49,
     RACK1, X49);

endmodule


// Library - XB16TSMC65, Cell - ZINVAI, View - schematic
// LAST TIME SAVED: May  8 15:13:02 2023
// NETLIST TIME: May 12 11:49:58 2023
`timescale 1ns / 1ns

module ZINVAI ( Z00, Z01, Z02, Z03, Z10, Z11, Z12, Z13, Z20, Z21, Z22,
     Z23, Z30, Z31, Z32, Z33, Z40, Z41, Z42, Z43, Z50, Z51, Z52, Z53,
     Z60, Z61, Z62, Z63, Z70, Z71, Z72, Z73, Z80, Z81, Z82, Z83, Z90,
     Z91, Z92, Z93, Z100, Z101, Z102, Z103, Z110, Z111, Z112, Z113,
     Z120, Z121, Z122, Z123, Z130, Z131, Z132, Z133, Z140, Z141, Z142,
     Z143, Z150, Z151, Z152, Z153, A00, A01, A02, A03, A10, A11, A12,
     A13, A20, A21, A22, A23, A30, A31, A32, A33, A40, A41, A42, A43,
     A50, A51, A52, A53, A60, A61, A62, A63, A70, A71, A72, A73, A80,
     A81, A82, A83, A90, A91, A92, A93, A100, A101, A102, A103, A110,
     A111, A112, A113, A120, A121, A122, A123, A130, A131, A132, A133,
     A140, A141, A142, A143, A150, A151, A152, A153 );

output  Z00, Z01, Z02, Z03, Z10, Z11, Z12, Z13, Z20, Z21, Z22, Z23,
     Z30, Z31, Z32, Z33, Z40, Z41, Z42, Z43, Z50, Z51, Z52, Z53, Z60,
     Z61, Z62, Z63, Z70, Z71, Z72, Z73, Z80, Z81, Z82, Z83, Z90, Z91,
     Z92, Z93, Z100, Z101, Z102, Z103, Z110, Z111, Z112, Z113, Z120,
     Z121, Z122, Z123, Z130, Z131, Z132, Z133, Z140, Z141, Z142, Z143,
     Z150, Z151, Z152, Z153;

input  A00, A01, A02, A03, A10, A11, A12, A13, A20, A21, A22, A23, A30,
     A31, A32, A33, A40, A41, A42, A43, A50, A51, A52, A53, A60, A61,
     A62, A63, A70, A71, A72, A73, A80, A81, A82, A83, A90, A91, A92,
     A93, A100, A101, A102, A103, A110, A111, A112, A113, A120, A121,
     A122, A123, A130, A131, A132, A133, A140, A141, A142, A143, A150,
     A151, A152, A153;


specify
    specparam CDS_LIBNAME  = "XB16TSMC65";
    specparam CDS_CELLNAME = "ZINVAI";
    specparam CDS_VIEWNAME = "schematic";
endspecify

INVXB1 I63 ( Z150, cds_globals.vdd_, cds_globals.gnd_, A150);
INVXB1 I62 ( Z151, cds_globals.vdd_, cds_globals.gnd_, A151);
INVXB1 I61 ( Z152, cds_globals.vdd_, cds_globals.gnd_, A152);
INVXB1 I60 ( Z153, cds_globals.vdd_, cds_globals.gnd_, A153);
INVXB1 I59 ( Z100, cds_globals.vdd_, cds_globals.gnd_, A100);
INVXB1 I58 ( Z101, cds_globals.vdd_, cds_globals.gnd_, A101);
INVXB1 I57 ( Z102, cds_globals.vdd_, cds_globals.gnd_, A102);
INVXB1 I56 ( Z103, cds_globals.vdd_, cds_globals.gnd_, A103);
INVXB1 I55 ( Z110, cds_globals.vdd_, cds_globals.gnd_, A110);
INVXB1 I54 ( Z111, cds_globals.vdd_, cds_globals.gnd_, A111);
INVXB1 I53 ( Z112, cds_globals.vdd_, cds_globals.gnd_, A112);
INVXB1 I52 ( Z113, cds_globals.vdd_, cds_globals.gnd_, A113);
INVXB1 I51 ( Z120, cds_globals.vdd_, cds_globals.gnd_, A120);
INVXB1 I50 ( Z121, cds_globals.vdd_, cds_globals.gnd_, A121);
INVXB1 I49 ( Z122, cds_globals.vdd_, cds_globals.gnd_, A122);
INVXB1 I48 ( Z123, cds_globals.vdd_, cds_globals.gnd_, A123);
INVXB1 I47 ( Z130, cds_globals.vdd_, cds_globals.gnd_, A130);
INVXB1 I46 ( Z131, cds_globals.vdd_, cds_globals.gnd_, A131);
INVXB1 I45 ( Z132, cds_globals.vdd_, cds_globals.gnd_, A132);
INVXB1 I44 ( Z133, cds_globals.vdd_, cds_globals.gnd_, A133);
INVXB1 I43 ( Z140, cds_globals.vdd_, cds_globals.gnd_, A140);
INVXB1 I42 ( Z141, cds_globals.vdd_, cds_globals.gnd_, A141);
INVXB1 I41 ( Z142, cds_globals.vdd_, cds_globals.gnd_, A142);
INVXB1 I40 ( Z143, cds_globals.vdd_, cds_globals.gnd_, A143);
INVXB1 I39 ( Z50, cds_globals.vdd_, cds_globals.gnd_, A50);
INVXB1 I38 ( Z51, cds_globals.vdd_, cds_globals.gnd_, A51);
INVXB1 I37 ( Z52, cds_globals.vdd_, cds_globals.gnd_, A52);
INVXB1 I36 ( Z53, cds_globals.vdd_, cds_globals.gnd_, A53);
INVXB1 I35 ( Z60, cds_globals.vdd_, cds_globals.gnd_, A60);
INVXB1 I34 ( Z61, cds_globals.vdd_, cds_globals.gnd_, A61);
INVXB1 I33 ( Z62, cds_globals.vdd_, cds_globals.gnd_, A62);
INVXB1 I32 ( Z63, cds_globals.vdd_, cds_globals.gnd_, A63);
INVXB1 I31 ( Z70, cds_globals.vdd_, cds_globals.gnd_, A70);
INVXB1 I30 ( Z71, cds_globals.vdd_, cds_globals.gnd_, A71);
INVXB1 I29 ( Z72, cds_globals.vdd_, cds_globals.gnd_, A72);
INVXB1 I28 ( Z73, cds_globals.vdd_, cds_globals.gnd_, A73);
INVXB1 I27 ( Z80, cds_globals.vdd_, cds_globals.gnd_, A80);
INVXB1 I26 ( Z81, cds_globals.vdd_, cds_globals.gnd_, A81);
INVXB1 I25 ( Z82, cds_globals.vdd_, cds_globals.gnd_, A82);
INVXB1 I24 ( Z83, cds_globals.vdd_, cds_globals.gnd_, A83);
INVXB1 I23 ( Z90, cds_globals.vdd_, cds_globals.gnd_, A90);
INVXB1 I22 ( Z91, cds_globals.vdd_, cds_globals.gnd_, A91);
INVXB1 I21 ( Z92, cds_globals.vdd_, cds_globals.gnd_, A92);
INVXB1 I20 ( Z93, cds_globals.vdd_, cds_globals.gnd_, A93);
INVXB1 I19 ( Z43, cds_globals.vdd_, cds_globals.gnd_, A43);
INVXB1 I18 ( Z42, cds_globals.vdd_, cds_globals.gnd_, A42);
INVXB1 I17 ( Z41, cds_globals.vdd_, cds_globals.gnd_, A41);
INVXB1 I16 ( Z40, cds_globals.vdd_, cds_globals.gnd_, A40);
INVXB1 I15 ( Z33, cds_globals.vdd_, cds_globals.gnd_, A33);
INVXB1 I14 ( Z32, cds_globals.vdd_, cds_globals.gnd_, A32);
INVXB1 I13 ( Z31, cds_globals.vdd_, cds_globals.gnd_, A31);
INVXB1 I12 ( Z30, cds_globals.vdd_, cds_globals.gnd_, A30);
INVXB1 I11 ( Z23, cds_globals.vdd_, cds_globals.gnd_, A23);
INVXB1 I10 ( Z22, cds_globals.vdd_, cds_globals.gnd_, A22);
INVXB1 I9 ( Z21, cds_globals.vdd_, cds_globals.gnd_, A21);
INVXB1 I8 ( Z20, cds_globals.vdd_, cds_globals.gnd_, A20);
INVXB1 I7 ( Z13, cds_globals.vdd_, cds_globals.gnd_, A13);
INVXB1 I6 ( Z12, cds_globals.vdd_, cds_globals.gnd_, A12);
INVXB1 I5 ( Z11, cds_globals.vdd_, cds_globals.gnd_, A11);
INVXB1 I4 ( Z10, cds_globals.vdd_, cds_globals.gnd_, A10);
INVXB1 I3 ( Z03, cds_globals.vdd_, cds_globals.gnd_, A03);
INVXB1 I2 ( Z02, cds_globals.vdd_, cds_globals.gnd_, A02);
INVXB1 I1 ( Z01, cds_globals.vdd_, cds_globals.gnd_, A01);
INVXB1 I0 ( Z00, cds_globals.vdd_, cds_globals.gnd_, A00);

endmodule


// Library - XB16TSMC65, Cell - ZLVL1R, View - schematic
// LAST TIME SAVED: May  8 15:13:02 2023
// NETLIST TIME: May 12 11:49:58 2023
`timescale 1ns / 1ns

module ZLVL1R ( Lval, L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11,
     L12, L13, L14, L15 );

output  Lval;

input  L0, L1, L2, L3, L4, L5, L6, L7, L8, L9, L10, L11, L12, L13, L14,
     L15;


specify
    specparam CDS_LIBNAME  = "XB16TSMC65";
    specparam CDS_CELLNAME = "ZLVL1R";
    specparam CDS_VIEWNAME = "schematic";
endspecify

INVXB1 I89 ( net014, cds_globals.vdd_, cds_globals.gnd_, net06);
INVXB1 I88 ( net013, cds_globals.vdd_, cds_globals.gnd_, net03);
INVXB1 I87 ( net04, cds_globals.vdd_, cds_globals.gnd_, net01);
INVXB1 I90 ( net012, cds_globals.vdd_, cds_globals.gnd_, net02);
INVXB1 I91 ( net026, cds_globals.vdd_, cds_globals.gnd_, net05);
ND4XB1 I81 ( net01, cds_globals.vdd_, cds_globals.gnd_, L0, L1, L2,
     L3);
ND4XB1 I82 ( net03, cds_globals.vdd_, cds_globals.gnd_, L4, L5, L6,
     L7);
ND4XB1 I85 ( net05, cds_globals.vdd_, cds_globals.gnd_, net022, net024,
     net025, net023);
ND4XB1 I84 ( net06, cds_globals.vdd_, cds_globals.gnd_, L8, L9, L10,
     L11);
ND4XB1 I83 ( net02, cds_globals.vdd_, cds_globals.gnd_, L12, L13, L14,
     L15);
INVXB2 I104 ( net07, cds_globals.vdd_, cds_globals.gnd_, net04);
INVXB2 I110 ( net010, cds_globals.vdd_, cds_globals.gnd_, net012);
INVXB2 I102 ( net020, cds_globals.vdd_, cds_globals.gnd_, net026);
INVXB2 I107 ( net08, cds_globals.vdd_, cds_globals.gnd_, net013);
INVXB2 I108 ( net09, cds_globals.vdd_, cds_globals.gnd_, net014);
INVXB4 I106 ( net024, cds_globals.vdd_, cds_globals.gnd_, net08);
INVXB4 I103 ( Lval, cds_globals.vdd_, cds_globals.gnd_, net020);
INVXB4 I105 ( net022, cds_globals.vdd_, cds_globals.gnd_, net07);
INVXB4 I111 ( net023, cds_globals.vdd_, cds_globals.gnd_, net010);
INVXB4 I109 ( net025, cds_globals.vdd_, cds_globals.gnd_, net09);

endmodule


// Library - XB16TSMC65, Cell - XB1616, View - schematic
// LAST TIME SAVED: May  9 14:24:20 2023
// NETLIST TIME: May 12 11:49:59 2023
`timescale 1ns / 1ns

module XB1616 ( LACK0, LACK1, LACK2, LACK3, LACK4, LACK5, LACK6, LACK7,
     LACK8, LACK9, LACK10, LACK11, LACK12, LACK13, LACK14, LACK15,
     LACKSE, NLACK0, NLACK1, NLACK2, NLACK3, NLACK4, NLACK5, NLACK6,
     NLACK7, NLACK8, NLACK9, NLACK10, NLACK11, NLACK12, NLACK13,
     NLACK14, NLACK15, NLACKSE, NR00, NR01, NR02, NR03, NR10, NR11,
     NR12, NR13, NR20, NR21, NR22, NR23, NR30, NR31, NR32, NR33, NR40,
     NR41, NR42, NR43, NR50, NR51, NR52, NR53, NR60, NR61, NR62, NR63,
     NR70, NR71, NR72, NR73, NR80, NR81, NR82, NR83, NR90, NR91, NR92,
     NR93, NR100, NR101, NR102, NR103, NR110, NR111, NR112, NR113,
     NR120, NR121, NR122, NR123, NR130, NR131, NR132, NR133, NR140,
     NR141, NR142, NR143, NR150, NR151, NR152, NR153, R00, R01, R02,
     R03, R10, R11, R12, R13, R20, R21, R22, R23, R30, R31, R32, R33,
     R40, R41, R42, R43, R50, R51, R52, R53, R60, R61, R62, R63, R70,
     R71, R72, R73, R80, R81, R82, R83, R90, R91, R92, R93, R100, R101,
     R102, R103, R110, R111, R112, R113, R120, R121, R122, R123, R130,
     R131, R132, R133, R140, R141, R142, R143, R150, R151, R152, R153,
     L00, L01, L02, L03, L10, L11, L12, L13, L20, L21, L22, L23, L30,
     L31, L32, L33, L40, L41, L42, L43, L50, L51, L52, L53, L60, L61,
     L62, L63, L70, L71, L72, L73, L80, L81, L82, L83, L90, L91, L92,
     L93, L100, L101, L102, L103, L110, L111, L112, L113, L120, L121,
     L122, L123, L130, L131, L132, L133, L140, L141, L142, L143, L150,
     L151, L152, L153, NL00, NL01, NL02, NL03, NL10, NL11, NL12, NL13,
     NL20, NL21, NL22, NL23, NL30, NL31, NL32, NL33, NL40, NL41, NL42,
     NL43, NL50, NL51, NL52, NL53, NL60, NL61, NL62, NL63, NL70, NL71,
     NL72, NL73, NL80, NL81, NL82, NL83, NL90, NL91, NL92, NL93, NL100,
     NL101, NL102, NL103, NL110, NL111, NL112, NL113, NL120, NL121,
     NL122, NL123, NL130, NL131, NL132, NL133, NL140, NL141, NL142,
     NL143, NL150, NL151, NL152, NL153, NRACK0, NRACK1, NRACK2, NRACK3,
     NRACK4, NRACK5, NRACK6, NRACK7, NRACK8, NRACK9, NRACK10, NRACK11,
     NRACK12, NRACK13, NRACK14, NRACK15, NX0, NX1, NX2, NX3, NX4, NX5,
     NX6, NX7, NX8, NX9, NX10, NX11, NX12, NX13, NX14, NX15, NX16,
     NX17, NX18, NX19, NX20, NX21, NX22, NX23, NX24, NX25, NX26, NX27,
     NX28, NX29, NX30, NX31, NX32, NX33, NX34, NX35, NX36, NX37, NX38,
     NX39, NX40, NX41, NX42, NX43, NX44, NX45, NX46, NX47, NX48, NX49,
     NX50, NX51, NX52, NX53, NX54, NX55, NX56, NX57, NX58, NX59, NX60,
     NX61, NX62, NX63, NX64, NX65, NX66, NX67, NX68, NX69, NX70, NX71,
     NX72, NX73, NX74, NX75, NX76, NX77, NX78, NX79, NX80, NX81, NX82,
     NX83, NX84, NX85, NX86, NX87, NX88, NX89, NX90, NX91, NX92, NX93,
     NX94, NX95, NX96, NX97, NX98, NX99, NX100, NX101, NX102, NX103,
     NX104, NX105, NX106, NX107, NX108, NX109, NX110, NX111, NX112,
     NX113, NX114, NX115, NX116, NX117, NX118, NX119, NX120, NX121,
     NX122, NX123, NX124, NX125, NX126, NX127, NX128, NX129, NX130,
     NX131, NX132, NX133, NX134, NX135, NX136, NX137, NX138, NX139,
     NX140, NX141, NX142, NX143, NX144, NX145, NX146, NX147, NX148,
     NX149, NX150, NX151, NX152, NX153, NX154, NX155, NX156, NX157,
     NX158, NX159, NX160, NX161, NX162, NX163, NX164, NX165, NX166,
     NX167, NX168, NX169, NX170, NX171, NX172, NX173, NX174, NX175,
     NX176, NX177, NX178, NX179, NX180, NX181, NX182, NX183, NX184,
     NX185, NX186, NX187, NX188, NX189, NX190, NX191, NX192, NX193,
     NX194, NX195, NX196, NX197, NX198, NX199, NX200, NX201, NX202,
     NX203, NX204, NX205, NX206, NX207, NX208, NX209, NX210, NX211,
     NX212, NX213, NX214, NX215, NX216, NX217, NX218, NX219, NX220,
     NX221, NX222, NX223, NX224, NX225, NX226, NX227, NX228, NX229,
     NX230, NX231, NX232, NX233, NX234, NX235, NX236, NX237, NX238,
     NX239, NX240, NX241, NX242, NX243, NX244, NX245, NX246, NX247,
     NX248, NX249, NX250, NX251, NX252, NX253, NX254, NX255, RACK0,
     RACK1, RACK2, RACK3, RACK4, RACK5, RACK6, RACK7, RACK8, RACK9,
     RACK10, RACK11, RACK12, RACK13, RACK14, RACK15, X0, X1, X2, X3,
     X4, X5, X6, X7, X8, X9, X10, X11, X12, X13, X14, X15, X16, X17,
     X18, X19, X20, X21, X22, X23, X24, X25, X26, X27, X28, X29, X30,
     X31, X32, X33, X34, X35, X36, X37, X38, X39, X40, X41, X42, X43,
     X44, X45, X46, X47, X48, X49, X50, X51, X52, X53, X54, X55, X56,
     X57, X58, X59, X60, X61, X62, X63, X64, X65, X66, X67, X68, X69,
     X70, X71, X72, X73, X74, X75, X76, X77, X78, X79, X80, X81, X82,
     X83, X84, X85, X86, X87, X88, X89, X90, X91, X92, X93, X94, X95,
     X96, X97, X98, X99, X100, X101, X102, X103, X104, X105, X106,
     X107, X108, X109, X110, X111, X112, X113, X114, X115, X116, X117,
     X118, X119, X120, X121, X122, X123, X124, X125, X126, X127, X128,
     X129, X130, X131, X132, X133, X134, X135, X136, X137, X138, X139,
     X140, X141, X142, X143, X144, X145, X146, X147, X148, X149, X150,
     X151, X152, X153, X154, X155, X156, X157, X158, X159, X160, X161,
     X162, X163, X164, X165, X166, X167, X168, X169, X170, X171, X172,
     X173, X174, X175, X176, X177, X178, X179, X180, X181, X182, X183,
     X184, X185, X186, X187, X188, X189, X190, X191, X192, X193, X194,
     X195, X196, X197, X198, X199, X200, X201, X202, X203, X204, X205,
     X206, X207, X208, X209, X210, X211, X212, X213, X214, X215, X216,
     X217, X218, X219, X220, X221, X222, X223, X224, X225, X226, X227,
     X228, X229, X230, X231, X232, X233, X234, X235, X236, X237, X238,
     X239, X240, X241, X242, X243, X244, X245, X246, X247, X248, X249,
     X250, X251, X252, X253, X254, X255 );

output  LACK0, LACK1, LACK2, LACK3, LACK4, LACK5, LACK6, LACK7, LACK8,
     LACK9, LACK10, LACK11, LACK12, LACK13, LACK14, LACK15, LACKSE,
     NLACK0, NLACK1, NLACK2, NLACK3, NLACK4, NLACK5, NLACK6, NLACK7,
     NLACK8, NLACK9, NLACK10, NLACK11, NLACK12, NLACK13, NLACK14,
     NLACK15, NLACKSE;

inout  NR00, NR01, NR02, NR03, NR10, NR11, NR12, NR13, NR20, NR21,
     NR22, NR23, NR30, NR31, NR32, NR33, NR40, NR41, NR42, NR43, NR50,
     NR51, NR52, NR53, NR60, NR61, NR62, NR63, NR70, NR71, NR72, NR73,
     NR80, NR81, NR82, NR83, NR90, NR91, NR92, NR93, NR100, NR101,
     NR102, NR103, NR110, NR111, NR112, NR113, NR120, NR121, NR122,
     NR123, NR130, NR131, NR132, NR133, NR140, NR141, NR142, NR143,
     NR150, NR151, NR152, NR153, R00, R01, R02, R03, R10, R11, R12,
     R13, R20, R21, R22, R23, R30, R31, R32, R33, R40, R41, R42, R43,
     R50, R51, R52, R53, R60, R61, R62, R63, R70, R71, R72, R73, R80,
     R81, R82, R83, R90, R91, R92, R93, R100, R101, R102, R103, R110,
     R111, R112, R113, R120, R121, R122, R123, R130, R131, R132, R133,
     R140, R141, R142, R143, R150, R151, R152, R153;

input  L00, L01, L02, L03, L10, L11, L12, L13, L20, L21, L22, L23, L30,
     L31, L32, L33, L40, L41, L42, L43, L50, L51, L52, L53, L60, L61,
     L62, L63, L70, L71, L72, L73, L80, L81, L82, L83, L90, L91, L92,
     L93, L100, L101, L102, L103, L110, L111, L112, L113, L120, L121,
     L122, L123, L130, L131, L132, L133, L140, L141, L142, L143, L150,
     L151, L152, L153, NL00, NL01, NL02, NL03, NL10, NL11, NL12, NL13,
     NL20, NL21, NL22, NL23, NL30, NL31, NL32, NL33, NL40, NL41, NL42,
     NL43, NL50, NL51, NL52, NL53, NL60, NL61, NL62, NL63, NL70, NL71,
     NL72, NL73, NL80, NL81, NL82, NL83, NL90, NL91, NL92, NL93, NL100,
     NL101, NL102, NL103, NL110, NL111, NL112, NL113, NL120, NL121,
     NL122, NL123, NL130, NL131, NL132, NL133, NL140, NL141, NL142,
     NL143, NL150, NL151, NL152, NL153, NRACK0, NRACK1, NRACK2, NRACK3,
     NRACK4, NRACK5, NRACK6, NRACK7, NRACK8, NRACK9, NRACK10, NRACK11,
     NRACK12, NRACK13, NRACK14, NRACK15, NX0, NX1, NX2, NX3, NX4, NX5,
     NX6, NX7, NX8, NX9, NX10, NX11, NX12, NX13, NX14, NX15, NX16,
     NX17, NX18, NX19, NX20, NX21, NX22, NX23, NX24, NX25, NX26, NX27,
     NX28, NX29, NX30, NX31, NX32, NX33, NX34, NX35, NX36, NX37, NX38,
     NX39, NX40, NX41, NX42, NX43, NX44, NX45, NX46, NX47, NX48, NX49,
     NX50, NX51, NX52, NX53, NX54, NX55, NX56, NX57, NX58, NX59, NX60,
     NX61, NX62, NX63, NX64, NX65, NX66, NX67, NX68, NX69, NX70, NX71,
     NX72, NX73, NX74, NX75, NX76, NX77, NX78, NX79, NX80, NX81, NX82,
     NX83, NX84, NX85, NX86, NX87, NX88, NX89, NX90, NX91, NX92, NX93,
     NX94, NX95, NX96, NX97, NX98, NX99, NX100, NX101, NX102, NX103,
     NX104, NX105, NX106, NX107, NX108, NX109, NX110, NX111, NX112,
     NX113, NX114, NX115, NX116, NX117, NX118, NX119, NX120, NX121,
     NX122, NX123, NX124, NX125, NX126, NX127, NX128, NX129, NX130,
     NX131, NX132, NX133, NX134, NX135, NX136, NX137, NX138, NX139,
     NX140, NX141, NX142, NX143, NX144, NX145, NX146, NX147, NX148,
     NX149, NX150, NX151, NX152, NX153, NX154, NX155, NX156, NX157,
     NX158, NX159, NX160, NX161, NX162, NX163, NX164, NX165, NX166,
     NX167, NX168, NX169, NX170, NX171, NX172, NX173, NX174, NX175,
     NX176, NX177, NX178, NX179, NX180, NX181, NX182, NX183, NX184,
     NX185, NX186, NX187, NX188, NX189, NX190, NX191, NX192, NX193,
     NX194, NX195, NX196, NX197, NX198, NX199, NX200, NX201, NX202,
     NX203, NX204, NX205, NX206, NX207, NX208, NX209, NX210, NX211,
     NX212, NX213, NX214, NX215, NX216, NX217, NX218, NX219, NX220,
     NX221, NX222, NX223, NX224, NX225, NX226, NX227, NX228, NX229,
     NX230, NX231, NX232, NX233, NX234, NX235, NX236, NX237, NX238,
     NX239, NX240, NX241, NX242, NX243, NX244, NX245, NX246, NX247,
     NX248, NX249, NX250, NX251, NX252, NX253, NX254, NX255, RACK0,
     RACK1, RACK2, RACK3, RACK4, RACK5, RACK6, RACK7, RACK8, RACK9,
     RACK10, RACK11, RACK12, RACK13, RACK14, RACK15, X0, X1, X2, X3,
     X4, X5, X6, X7, X8, X9, X10, X11, X12, X13, X14, X15, X16, X17,
     X18, X19, X20, X21, X22, X23, X24, X25, X26, X27, X28, X29, X30,
     X31, X32, X33, X34, X35, X36, X37, X38, X39, X40, X41, X42, X43,
     X44, X45, X46, X47, X48, X49, X50, X51, X52, X53, X54, X55, X56,
     X57, X58, X59, X60, X61, X62, X63, X64, X65, X66, X67, X68, X69,
     X70, X71, X72, X73, X74, X75, X76, X77, X78, X79, X80, X81, X82,
     X83, X84, X85, X86, X87, X88, X89, X90, X91, X92, X93, X94, X95,
     X96, X97, X98, X99, X100, X101, X102, X103, X104, X105, X106,
     X107, X108, X109, X110, X111, X112, X113, X114, X115, X116, X117,
     X118, X119, X120, X121, X122, X123, X124, X125, X126, X127, X128,
     X129, X130, X131, X132, X133, X134, X135, X136, X137, X138, X139,
     X140, X141, X142, X143, X144, X145, X146, X147, X148, X149, X150,
     X151, X152, X153, X154, X155, X156, X157, X158, X159, X160, X161,
     X162, X163, X164, X165, X166, X167, X168, X169, X170, X171, X172,
     X173, X174, X175, X176, X177, X178, X179, X180, X181, X182, X183,
     X184, X185, X186, X187, X188, X189, X190, X191, X192, X193, X194,
     X195, X196, X197, X198, X199, X200, X201, X202, X203, X204, X205,
     X206, X207, X208, X209, X210, X211, X212, X213, X214, X215, X216,
     X217, X218, X219, X220, X221, X222, X223, X224, X225, X226, X227,
     X228, X229, X230, X231, X232, X233, X234, X235, X236, X237, X238,
     X239, X240, X241, X242, X243, X244, X245, X246, X247, X248, X249,
     X250, X251, X252, X253, X254, X255;


specify
    specparam CDS_LIBNAME  = "XB16TSMC65";
    specparam CDS_CELLNAME = "XB1616";
    specparam CDS_VIEWNAME = "schematic";
endspecify

ZLVL1R I27 ( LVAL3, NL03, NL13, NL23, NL33, NL43, NL53, NL63, NL73,
     NL83, NL93, NL103, NL113, NL123, NL133, NL143, NL153);
ZLVL1R I26 ( LVAL2, NL02, NL12, NL22, NL32, NL42, NL52, NL62, NL72,
     NL82, NL92, NL102, NL112, NL122, NL132, NL142, NL152);
ZLVL1R I25 ( LVAL1, NL01, NL11, NL21, NL31, NL41, NL51, NL61, NL71,
     NL81, NL91, NL101, NL111, NL121, NL131, NL141, NL151);
ZLVL1R I24 ( LVAL0, NL00, NL10, NL20, NL30, NL40, NL50, NL60, NL70,
     NL80, NL90, NL100, NL110, NL120, NL130, NL140, NL150);
ZRVLAR I44 ( net842, R00, R01, R02, R03, R10, R11, R12, R13, R20, R21,
     R22, R23, R30, R31, R32, R33, R40, R41, R42, R43, R50, R51, R52,
     R53, R60, R61, R62, R63, R70, R71, R72, R73, R80, R81, R82, R83,
     R90, R91, R92, R93, R100, R101, R102, R103, R110, R111, R112,
     R113, R120, R121, R122, R123, R130, R131, R132, R133, R140, R141,
     R142, R143, R150, R151, R152, R153);
ZFBAR4 I22 ( NR00, NR01, NR02, NR03, NR10, NR11, NR12, NR13, NR20,
     NR21, NR22, NR23, NR30, NR31, NR32, NR33, NR40, NR41, NR42, NR43,
     NR50, NR51, NR52, NR53, NR60, NR61, NR62, NR63, NR70, NR71, NR72,
     NR73, NR80, NR81, NR82, NR83, NR90, NR91, NR92, NR93, NR100,
     NR101, NR102, NR103, NR110, NR111, NR112, NR113, NR120, NR121,
     NR122, NR123, NR130, NR131, NR132, NR133, NR140, NR141, NR142,
     NR143, NR150, NR151, NR152, NR153, R00, R01, R02, R03, R10, R11,
     R12, R13, R20, R21, R22, R23, R30, R31, R32, R33, R40, R41, R42,
     R43, R50, R51, R52, R53, R60, R61, R62, R63, R70, R71, R72, R73,
     R80, R81, R82, R83, R90, R91, R92, R93, R100, R101, R102, R103,
     R110, R111, R112, R113, R120, R121, R122, R123, R130, R131, R132,
     R133, R140, R141, R142, R143, R150, R151, R152, R153,
     cds_globals.vdda_, cds_globals.gnd_, L00, L01, L02, L03, L10, L11,
     L12, L13, L20, L21, L22, L23, L30, L31, L32, L33, L40, L41, L42,
     L43, L50, L51, L52, L53, L60, L61, L62, L63, L70, L71, L72, L73,
     L80, L81, L82, L83, L90, L91, L92, L93, L100, L101, L102, L103,
     L110, L111, L112, L113, L120, L121, L122, L123, L130, L131, L132,
     L133, L140, L141, L142, L143, L150, L151, L152, L153, NL00, NL01,
     NL02, NL03, NL10, NL11, NL12, NL13, NL20, NL21, NL22, NL23, NL30,
     NL31, NL32, NL33, NL40, NL41, NL42, NL43, NL50, NL51, NL52, NL53,
     NL60, NL61, NL62, NL63, NL70, NL71, NL72, NL73, NL80, NL81, NL82,
     NL83, NL90, NL91, NL92, NL93, NL100, NL101, NL102, NL103, NL110,
     NL111, NL112, NL113, NL120, NL121, NL122, NL123, NL130, NL131,
     NL132, NL133, NL140, NL141, NL142, NL143, NL150, NL151, NL152,
     NL153, NRACK0, NRACK1, NRACK2, NRACK3, NRACK4, NRACK5, NRACK6,
     NRACK7, NRACK8, NRACK9, NRACK10, NRACK11, NRACK12, NRACK13,
     NRACK14, NRACK15, LVAL0, LVAL1, LVAL2, LVAL3, NX0, NX1, NX2, NX3,
     NX4, NX5, NX6, NX7, NX8, NX9, NX10, NX11, NX12, NX13, NX14, NX15,
     NX16, NX17, NX18, NX19, NX20, NX21, NX22, NX23, NX24, NX25, NX26,
     NX27, NX28, NX29, NX30, NX31, NX32, NX33, NX34, NX35, NX36, NX37,
     NX38, NX39, NX40, NX41, NX42, NX43, NX44, NX45, NX46, NX47, NX48,
     NX49, NX50, NX51, NX52, NX53, NX54, NX55, NX56, NX57, NX58, NX59,
     NX60, NX61, NX62, NX63, NX64, NX65, NX66, NX67, NX68, NX69, NX70,
     NX71, NX72, NX73, NX74, NX75, NX76, NX77, NX78, NX79, NX80, NX81,
     NX82, NX83, NX84, NX85, NX86, NX87, NX88, NX89, NX90, NX91, NX92,
     NX93, NX94, NX95, NX96, NX97, NX98, NX99, NX100, NX101, NX102,
     NX103, NX104, NX105, NX106, NX107, NX108, NX109, NX110, NX111,
     NX112, NX113, NX114, NX115, NX116, NX117, NX118, NX119, NX120,
     NX121, NX122, NX123, NX124, NX125, NX126, NX127, NX128, NX129,
     NX130, NX131, NX132, NX133, NX134, NX135, NX136, NX137, NX138,
     NX139, NX140, NX141, NX142, NX143, NX144, NX145, NX146, NX147,
     NX148, NX149, NX150, NX151, NX152, NX153, NX154, NX155, NX156,
     NX157, NX158, NX159, NX160, NX161, NX162, NX163, NX164, NX165,
     NX166, NX167, NX168, NX169, NX170, NX171, NX172, NX173, NX174,
     NX175, NX176, NX177, NX178, NX179, NX180, NX181, NX182, NX183,
     NX184, NX185, NX186, NX187, NX188, NX189, NX190, NX191, NX192,
     NX193, NX194, NX195, NX196, NX197, NX198, NX199, NX200, NX201,
     NX202, NX203, NX204, NX205, NX206, NX207, NX208, NX209, NX210,
     NX211, NX212, NX213, NX214, NX215, NX216, NX217, NX218, NX219,
     NX220, NX221, NX222, NX223, NX224, NX225, NX226, NX227, NX228,
     NX229, NX230, NX231, NX232, NX233, NX234, NX235, NX236, NX237,
     NX238, NX239, NX240, NX241, NX242, NX243, NX244, NX245, NX246,
     NX247, NX248, NX249, NX250, NX251, NX252, NX253, NX254, NX255,
     RACK0, RACK1, RACK2, RACK3, RACK4, RACK5, RACK6, RACK7, RACK8,
     RACK9, RACK10, RACK11, RACK12, RACK13, RACK14, RACK15, X0, X1, X2,
     X3, X4, X5, X6, X7, X8, X9, X10, X11, X12, X13, X14, X15, X16,
     X17, X18, X19, X20, X21, X22, X23, X24, X25, X26, X27, X28, X29,
     X30, X31, X32, X33, X34, X35, X36, X37, X38, X39, X40, X41, X42,
     X43, X44, X45, X46, X47, X48, X49, X50, X51, X52, X53, X54, X55,
     X56, X57, X58, X59, X60, X61, X62, X63, X64, X65, X66, X67, X68,
     X69, X70, X71, X72, X73, X74, X75, X76, X77, X78, X79, X80, X81,
     X82, X83, X84, X85, X86, X87, X88, X89, X90, X91, X92, X93, X94,
     X95, X96, X97, X98, X99, X100, X101, X102, X103, X104, X105, X106,
     X107, X108, X109, X110, X111, X112, X113, X114, X115, X116, X117,
     X118, X119, X120, X121, X122, X123, X124, X125, X126, X127, X128,
     X129, X130, X131, X132, X133, X134, X135, X136, X137, X138, X139,
     X140, X141, X142, X143, X144, X145, X146, X147, X148, X149, X150,
     X151, X152, X153, X154, X155, X156, X157, X158, X159, X160, X161,
     X162, X163, X164, X165, X166, X167, X168, X169, X170, X171, X172,
     X173, X174, X175, X176, X177, X178, X179, X180, X181, X182, X183,
     X184, X185, X186, X187, X188, X189, X190, X191, X192, X193, X194,
     X195, X196, X197, X198, X199, X200, X201, X202, X203, X204, X205,
     X206, X207, X208, X209, X210, X211, X212, X213, X214, X215, X216,
     X217, X218, X219, X220, X221, X222, X223, X224, X225, X226, X227,
     X228, X229, X230, X231, X232, X233, X234, X235, X236, X237, X238,
     X239, X240, X241, X242, X243, X244, X245, X246, X247, X248, X249,
     X250, X251, X252, X253, X254, X255);
ZINVAI I47 ( NR00, NR01, NR02, NR03, NR10, NR11, NR12, NR13, NR20,
     NR21, NR22, NR23, NR30, NR31, NR32, NR33, NR40, NR41, NR42, NR43,
     NR50, NR51, NR52, NR53, NR60, NR61, NR62, NR63, NR70, NR71, NR72,
     NR73, NR80, NR81, NR82, NR83, NR90, NR91, NR92, NR93, NR100,
     NR101, NR102, NR113, NR110, NR111, NR112, NR113, NR120, NR121,
     NR122, NR123, NR130, NR131, NR132, NR133, NR140, NR141, NR142,
     NR143, NR150, NR151, NR152, NR153, R00, R01, R02, R03, R10, R11,
     R12, R13, R20, R21, R22, R23, R30, R31, R32, R33, R40, R41, R42,
     R43, R50, R51, R52, R53, R60, R61, R62, R63, R70, R71, R72, R73,
     R80, R81, R82, R83, R90, R91, R92, R93, R100, R101, R102, R103,
     R110, R111, R112, R113, R120, R121, R122, R123, R130, R131, R132,
     R133, R140, R141, R142, R143, R150, R151, R152, R153);
ZLCKAO I45 ( LACK0, LACK1, LACK2, LACK3, LACK4, LACK5, LACK6, LACK7,
     LACK8, LACK9, LACK10, LACK11, LACK12, LACK13, LACK14, LACK15, E0,
     E1, E2, E3, E4, E5, E6, E7, E8, E9, E10, E11, E12, E13, E14, E15,
     net842);
ZCLAR4 I23 ( NR00, NR01, NR02, NR03, NR10, NR11, NR12, NR13, NR20,
     NR21, NR22, NR23, NR30, NR31, NR32, NR33, NR40, NR41, NR42, NR43,
     NR50, NR51, NR52, NR53, NR60, NR61, NR62, NR63, NR70, NR71, NR72,
     NR73, NR80, NR81, NR82, NR83, NR90, NR91, NR92, NR93, NR100,
     NR101, NR102, NR103, NR110, NR111, NR112, NR113, NR120, NR121,
     NR122, NR123, NR130, NR131, NR132, NR133, NR140, NR141, NR142,
     NR143, NR150, NR151, NR152, NR153, R00, R01, R02, R03, R10, R11,
     R12, R13, R20, R21, R22, R23, R30, R31, R32, R33, R40, R41, R42,
     R43, R50, R51, R52, R53, R60, R61, R62, R63, R70, R71, R72, R73,
     R80, R81, R82, R83, R90, R91, R92, R93, R100, R101, R102, R103,
     R110, R111, R112, R113, R120, R121, R122, R123, R130, R131, R132,
     R133, R140, R141, R142, R143, R150, R151, R152, R153,
     cds_globals.vdd_, cds_globals.gnd_, LVAL0, LVAL1, LVAL2, LVAL3,
     RACK0, RACK1, RACK2, RACK3, RACK4, RACK5, RACK6, RACK7, RACK8,
     RACK9, RACK10, RACK11, RACK12, RACK13, RACK14, RACK15);
ZXGNAX I46 ( E0, E1, E2, E3, E4, E5, E6, E7, E8, E9, E10, E11, E12,
     E13, E14, E15, X0, X1, X2, X3, X4, X5, X6, X7, X8, X9, X10, X11,
     X12, X13, X14, X15, X16, X17, X18, X19, X20, X21, X22, X23, X24,
     X25, X26, X27, X28, X29, X30, X31, X32, X33, X34, X35, X36, X37,
     X38, X39, X40, X41, X42, X43, X44, X45, X46, X47, X48, X49, X50,
     X51, X52, X53, X54, X55, X56, X57, X58, X59, X60, X61, X62, X63,
     X64, X65, X66, X67, X68, X69, X70, X71, X72, X73, X74, X75, X76,
     X77, X78, X79, X80, X81, X82, X83, X84, X85, X86, X87, X88, X89,
     X90, X91, X92, X93, X94, X95, X96, X97, X98, X99, X100, X101,
     X102, X103, X104, X105, X106, X107, X108, X109, X110, X111, X112,
     X113, X114, X115, X116, X117, X118, X119, X120, X121, X122, X123,
     X124, X125, X126, X127, X128, X129, X130, X131, X132, X133, X134,
     X135, X136, X137, X138, X139, X140, X141, X142, X143, X144, X145,
     X146, X147, X148, X149, X150, X151, X152, X153, X154, X155, X156,
     X157, X158, X159, X160, X161, X162, X163, X164, X165, X166, X167,
     X168, X169, X170, X171, X172, X173, X174, X175, X176, X177, X178,
     X179, X180, X181, X182, X183, X184, X185, X186, X187, X188, X189,
     X190, X191, X192, X193, X194, X195, X196, X197, X198, X199, X200,
     X201, X202, X203, X204, X205, X206, X207, X208, X209, X210, X211,
     X212, X213, X214, X215, X216, X217, X218, X219, X220, X221, X222,
     X223, X224, X225, X226, X227, X228, X229, X230, X231, X232, X233,
     X234, X235, X236, X237, X238, X239, X240, X241, X242, X243, X244,
     X245, X246, X247, X248, X249, X250, X251, X252, X253, X254, X255);

endmodule
